// Copyright 2022 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Fabian Schuiki <fschuiki@iis.ee.ethz.ch>
// Florian Zaruba <zarubaf@iis.ee.ethz.ch>
// Stefan Mach <smach@iis.ee.ethz.ch>
// Thomas Benz <tbenz@iis.ee.ethz.ch>
// Paul Scheffler <paulsc@iis.ee.ethz.ch>
// Wolfgang Roenninger <wroennin@iis.ee.ethz.ch>
//
// AUTOMATICALLY GENERATED by gen_bootrom.py; edit the script instead.

module cheshire_bootrom #(
    parameter int unsigned AddrWidth = 32,
    parameter int unsigned DataWidth = 32
)(
    input  logic                 clk_i,
    input  logic                 rst_ni,
    input  logic                 req_i,
    input  logic [AddrWidth-1:0] addr_i,
    output logic [DataWidth-1:0] data_o
);
    localparam unsigned NumWords = 4096;
    logic [$clog2(NumWords)-1:0] word;

    assign word = addr_i / (DataWidth / 8);

    always_comb begin
        data_o = '0;
        unique case (word)
        000: data_o = 32'h6f006117 /* 0x0000 */;
            001: data_o = 32'h00010113 /* 0x0004 */;
            002: data_o = 32'h00002197 /* 0x0008 */;
            003: data_o = 32'h39418193 /* 0x000c */;
            004: data_o = 32'h301012f3 /* 0x0010 */;
            005: data_o = 32'h0282f313 /* 0x0014 */;
            006: data_o = 32'h0082f293 /* 0x0018 */;
            007: data_o = 32'hfd830313 /* 0x001c */;
            008: data_o = 32'h0e031863 /* 0x0020 */;
            009: data_o = 32'h03364305 /* 0x0024 */;
            010: data_o = 32'h30032073 /* 0x0028 */;
            011: data_o = 32'hd2207053 /* 0x002c */;
            012: data_o = 32'hd22070d3 /* 0x0030 */;
            013: data_o = 32'hd2207153 /* 0x0034 */;
            014: data_o = 32'hd22071d3 /* 0x0038 */;
            015: data_o = 32'hd2207253 /* 0x003c */;
            016: data_o = 32'hd22072d3 /* 0x0040 */;
            017: data_o = 32'hd2207353 /* 0x0044 */;
            018: data_o = 32'hd22073d3 /* 0x0048 */;
            019: data_o = 32'hd2207453 /* 0x004c */;
            020: data_o = 32'hd22074d3 /* 0x0050 */;
            021: data_o = 32'hd2207553 /* 0x0054 */;
            022: data_o = 32'hd22075d3 /* 0x0058 */;
            023: data_o = 32'hd2207653 /* 0x005c */;
            024: data_o = 32'hd22076d3 /* 0x0060 */;
            025: data_o = 32'hd2207753 /* 0x0064 */;
            026: data_o = 32'hd22077d3 /* 0x0068 */;
            027: data_o = 32'hd2207853 /* 0x006c */;
            028: data_o = 32'hd22078d3 /* 0x0070 */;
            029: data_o = 32'hd2207953 /* 0x0074 */;
            030: data_o = 32'hd22079d3 /* 0x0078 */;
            031: data_o = 32'hd2207a53 /* 0x007c */;
            032: data_o = 32'hd2207ad3 /* 0x0080 */;
            033: data_o = 32'hd2207b53 /* 0x0084 */;
            034: data_o = 32'hd2207bd3 /* 0x0088 */;
            035: data_o = 32'hd2207c53 /* 0x008c */;
            036: data_o = 32'hd2207cd3 /* 0x0090 */;
            037: data_o = 32'hd2207d53 /* 0x0094 */;
            038: data_o = 32'hd2207dd3 /* 0x0098 */;
            039: data_o = 32'hd2207e53 /* 0x009c */;
            040: data_o = 32'hd2207ed3 /* 0x00a0 */;
            041: data_o = 32'hd2207f53 /* 0x00a4 */;
            042: data_o = 32'hd2207fd3 /* 0x00a8 */;
            043: data_o = 32'h30033073 /* 0x00ac */;
            044: data_o = 32'h42014081 /* 0x00b0 */;
            045: data_o = 32'h43014281 /* 0x00b4 */;
            046: data_o = 32'h44014381 /* 0x00b8 */;
            047: data_o = 32'h45014481 /* 0x00bc */;
            048: data_o = 32'h46014581 /* 0x00c0 */;
            049: data_o = 32'h47014681 /* 0x00c4 */;
            050: data_o = 32'h48014781 /* 0x00c8 */;
            051: data_o = 32'h49014881 /* 0x00cc */;
            052: data_o = 32'h4a014981 /* 0x00d0 */;
            053: data_o = 32'h4b014a81 /* 0x00d4 */;
            054: data_o = 32'h4c014b81 /* 0x00d8 */;
            055: data_o = 32'h4d014c81 /* 0x00dc */;
            056: data_o = 32'h4e014d81 /* 0x00e0 */;
            057: data_o = 32'h4f014e81 /* 0x00e4 */;
            058: data_o = 32'h12974f81 /* 0x00e8 */;
            059: data_o = 32'h82930100 /* 0x00ec */;
            060: data_o = 32'h537df162 /* 0x00f0 */;
            061: data_o = 32'h0062a023 /* 0x00f4 */;
            062: data_o = 32'h0062a223 /* 0x00f8 */;
            063: data_o = 32'ha8234305 /* 0x00fc */;
            064: data_o = 32'h42810062 /* 0x0100 */;
            065: data_o = 32'h100f4301 /* 0x0104 */;
            066: data_o = 32'h10ef0000 /* 0x0108 */;
            067: data_o = 32'ha8514ef0 /* 0x010c */;
            068: data_o = 32'hfa0280e3 /* 0x0110 */;
            069: data_o = 32'h03364305 /* 0x0114 */;
            070: data_o = 32'h30032073 /* 0x0118 */;
            071: data_o = 32'hd0207053 /* 0x011c */;
            072: data_o = 32'hd02070d3 /* 0x0120 */;
            073: data_o = 32'hd0207153 /* 0x0124 */;
            074: data_o = 32'hd02071d3 /* 0x0128 */;
            075: data_o = 32'hd0207253 /* 0x012c */;
            076: data_o = 32'hd02072d3 /* 0x0130 */;
            077: data_o = 32'hd0207353 /* 0x0134 */;
            078: data_o = 32'hd02073d3 /* 0x0138 */;
            079: data_o = 32'hd0207453 /* 0x013c */;
            080: data_o = 32'hd02074d3 /* 0x0140 */;
            081: data_o = 32'hd0207553 /* 0x0144 */;
            082: data_o = 32'hd02075d3 /* 0x0148 */;
            083: data_o = 32'hd0207653 /* 0x014c */;
            084: data_o = 32'hd02076d3 /* 0x0150 */;
            085: data_o = 32'hd0207753 /* 0x0154 */;
            086: data_o = 32'hd02077d3 /* 0x0158 */;
            087: data_o = 32'hd0207853 /* 0x015c */;
            088: data_o = 32'hd02078d3 /* 0x0160 */;
            089: data_o = 32'hd0207953 /* 0x0164 */;
            090: data_o = 32'hd02079d3 /* 0x0168 */;
            091: data_o = 32'hd0207a53 /* 0x016c */;
            092: data_o = 32'hd0207ad3 /* 0x0170 */;
            093: data_o = 32'hd0207b53 /* 0x0174 */;
            094: data_o = 32'hd0207bd3 /* 0x0178 */;
            095: data_o = 32'hd0207c53 /* 0x017c */;
            096: data_o = 32'hd0207cd3 /* 0x0180 */;
            097: data_o = 32'hd0207d53 /* 0x0184 */;
            098: data_o = 32'hd0207dd3 /* 0x0188 */;
            099: data_o = 32'hd0207e53 /* 0x018c */;
            100: data_o = 32'hd0207ed3 /* 0x0190 */;
            101: data_o = 32'hd0207f53 /* 0x0194 */;
            102: data_o = 32'hd0207fd3 /* 0x0198 */;
            103: data_o = 32'h30033073 /* 0x019c */;
            104: data_o = 32'h0506bf01 /* 0x01a0 */;
            105: data_o = 32'h00156513 /* 0x01a4 */;
            106: data_o = 32'h01000297 /* 0x01a8 */;
            107: data_o = 32'he5828293 /* 0x01ac */;
            108: data_o = 32'h00a2a223 /* 0x01b0 */;
            109: data_o = 32'h10500073 /* 0x01b4 */;
            110: data_o = 32'h832abff5 /* 0x01b8 */;
            111: data_o = 32'h0023c611 /* 0x01bc */;
            112: data_o = 32'h167d00b3 /* 0x01c0 */;
            113: data_o = 32'hfe650305 /* 0x01c4 */;
            114: data_o = 32'hc9098082 /* 0x01c8 */;
            115: data_o = 32'h4501611c /* 0x01cc */;
            116: data_o = 32'h27814f9c /* 0x01d0 */;
            117: data_o = 32'h8023c589 /* 0x01d4 */;
            118: data_o = 32'h808200f5 /* 0x01d8 */;
            119: data_o = 32'h80824509 /* 0x01dc */;
            120: data_o = 32'h3797cd11 /* 0x01e0 */;
            121: data_o = 32'h87930100 /* 0x01e4 */;
            122: data_o = 32'hc783e1e7 /* 0x01e8 */;
            123: data_o = 32'hf7930147 /* 0x01ec */;
            124: data_o = 32'hdbe50207 /* 0x01f0 */;
            125: data_o = 32'h01003797 /* 0x01f4 */;
            126: data_o = 32'he0a78623 /* 0x01f8 */;
            127: data_o = 32'h78138082 /* 0x01fc */;
            128: data_o = 32'h47810026 /* 0x0200 */;
            129: data_o = 32'h17638a05 /* 0x0204 */;
            130: data_o = 32'h49580008 /* 0x0208 */;
            131: data_o = 32'he3194785 /* 0x020c */;
            132: data_o = 32'h0006079b /* 0x0210 */;
            133: data_o = 32'h4705c611 /* 0x0214 */;
            134: data_o = 32'h4914c958 /* 0x0218 */;
            135: data_o = 32'hd3146118 /* 0x021c */;
            136: data_o = 32'h1463e595 /* 0x0220 */;
            137: data_o = 32'h45010008 /* 0x0224 */;
            138: data_o = 32'h491c8082 /* 0x0228 */;
            139: data_o = 32'h61181141 /* 0x022c */;
            140: data_o = 32'h2785e406 /* 0x0230 */;
            141: data_o = 32'h00052a23 /* 0x0234 */;
            142: data_o = 32'hd31c8b85 /* 0x0238 */;
            143: data_o = 32'h45a14601 /* 0x023c */;
            144: data_o = 32'hfbfff0ef /* 0x0240 */;
            145: data_o = 32'h450160a2 /* 0x0244 */;
            146: data_o = 32'h80820141 /* 0x0248 */;
            147: data_o = 32'h67096114 /* 0x024c */;
            148: data_o = 32'h71070713 /* 0x0250 */;
            149: data_o = 32'h46634ad0 /* 0x0254 */;
            150: data_o = 32'h377d0006 /* 0x0258 */;
            151: data_o = 32'h557dff65 /* 0x025c */;
            152: data_o = 32'hf5938082 /* 0x0260 */;
            153: data_o = 32'h35fd1ff5 /* 0x0264 */;
            154: data_o = 32'h0097979b /* 0x0268 */;
            155: data_o = 32'h25818ddd /* 0x026c */;
            156: data_o = 32'h0737d2cc /* 0x0270 */;
            157: data_o = 32'h4adc4000 /* 0x0274 */;
            158: data_o = 32'h27818ff9 /* 0x0278 */;
            159: data_o = 32'h04e3ffed /* 0x027c */;
            160: data_o = 32'h491cfa08 /* 0x0280 */;
            161: data_o = 32'h00052a23 /* 0x0284 */;
            162: data_o = 32'h8b852785 /* 0x0288 */;
            163: data_o = 32'hbf61d29c /* 0x028c */;
            164: data_o = 32'h882a87b2 /* 0x0290 */;
            165: data_o = 32'h863a8e2e /* 0x0294 */;
            166: data_o = 32'he291e399 /* 0x0298 */;
            167: data_o = 32'h7513b78d /* 0x029c */;
            168: data_o = 32'hc119007e /* 0x02a0 */;
            169: data_o = 32'h8082557d /* 0x02a4 */;
            170: data_o = 32'h78937179 /* 0x02a8 */;
            171: data_o = 32'hf4060026 /* 0x02ac */;
            172: data_o = 32'hec26f022 /* 0x02b0 */;
            173: data_o = 32'h4f018a05 /* 0x02b4 */;
            174: data_o = 32'h00089863 /* 0x02b8 */;
            175: data_o = 32'h01482703 /* 0x02bc */;
            176: data_o = 32'he3194f05 /* 0x02c0 */;
            177: data_o = 32'h00060f1b /* 0x02c4 */;
            178: data_o = 32'h4705ca09 /* 0x02c8 */;
            179: data_o = 32'h00e82a23 /* 0x02cc */;
            180: data_o = 32'h01082603 /* 0x02d0 */;
            181: data_o = 32'h00083703 /* 0x02d4 */;
            182: data_o = 32'h1563d310 /* 0x02d8 */;
            183: data_o = 32'h9463020e /* 0x02dc */;
            184: data_o = 32'h45010008 /* 0x02e0 */;
            185: data_o = 32'h2783a8d1 /* 0x02e4 */;
            186: data_o = 32'h37030108 /* 0x02e8 */;
            187: data_o = 32'h2a230008 /* 0x02ec */;
            188: data_o = 32'h27850008 /* 0x02f0 */;
            189: data_o = 32'hd31c8b85 /* 0x02f4 */;
            190: data_o = 32'h45a14601 /* 0x02f8 */;
            191: data_o = 32'hf0ef8542 /* 0x02fc */;
            192: data_o = 32'hb7c5f01f /* 0x0300 */;
            193: data_o = 32'h00f03733 /* 0x0304 */;
            194: data_o = 32'h0017171b /* 0x0308 */;
            195: data_o = 32'h00d03633 /* 0x030c */;
            196: data_o = 32'h1e9b8f51 /* 0x0310 */;
            197: data_o = 32'h571b0187 /* 0x0314 */;
            198: data_o = 32'h77130017 /* 0x0318 */;
            199: data_o = 32'h531b0ff7 /* 0x031c */;
            200: data_o = 32'h559b003e /* 0x0320 */;
            201: data_o = 32'hde9b003e /* 0x0324 */;
            202: data_o = 32'h3e03418e /* 0x0328 */;
            203: data_o = 32'hcf390008 /* 0x032c */;
            204: data_o = 32'h4023529b /* 0x0330 */;
            205: data_o = 32'h873e8616 /* 0x0334 */;
            206: data_o = 32'hf3934f81 /* 0x0338 */;
            207: data_o = 32'hf4130037 /* 0x033c */;
            208: data_o = 32'h90630017 /* 0x0340 */;
            209: data_o = 32'h1f9b09f2 /* 0x0344 */;
            210: data_o = 32'h877e0026 /* 0x0348 */;
            211: data_o = 32'h04bfd063 /* 0x034c */;
            212: data_o = 32'h01884603 /* 0x0350 */;
            213: data_o = 32'hcf8397fe /* 0x0354 */;
            214: data_o = 32'h073b0007 /* 0x0358 */;
            215: data_o = 32'hea7940e3 /* 0x035c */;
            216: data_o = 32'h01f105a3 /* 0x0360 */;
            217: data_o = 32'h4f814285 /* 0x0364 */;
            218: data_o = 32'h00e2d463 /* 0x0368 */;
            219: data_o = 32'h0017cf83 /* 0x036c */;
            220: data_o = 32'h01f10523 /* 0x0370 */;
            221: data_o = 32'h14634f8d /* 0x0374 */;
            222: data_o = 32'hc60301f7 /* 0x0378 */;
            223: data_o = 32'h04a30027 /* 0x037c */;
            224: data_o = 32'h042300c1 /* 0x0380 */;
            225: data_o = 32'h47a20001 /* 0x0384 */;
            226: data_o = 32'h02fe2423 /* 0x0388 */;
            227: data_o = 32'hfff3079b /* 0x038c */;
            228: data_o = 32'h00ce971b /* 0x0390 */;
            229: data_o = 32'h1ff7f793 /* 0x0394 */;
            230: data_o = 32'h1f1b8fd9 /* 0x0398 */;
            231: data_o = 32'he7b3009f /* 0x039c */;
            232: data_o = 32'h670901e7 /* 0x03a0 */;
            233: data_o = 32'h07132781 /* 0x03a4 */;
            234: data_o = 32'h26037107 /* 0x03a8 */;
            235: data_o = 32'h4363014e /* 0x03ac */;
            236: data_o = 32'h377d2006 /* 0x03b0 */;
            237: data_o = 32'h557dfb7d /* 0x03b4 */;
            238: data_o = 32'h740270a2 /* 0x03b8 */;
            239: data_o = 32'h614564e2 /* 0x03bc */;
            240: data_o = 32'h44838082 /* 0x03c0 */;
            241: data_o = 32'he49d0188 /* 0x03c4 */;
            242: data_o = 32'h00074483 /* 0x03c8 */;
            243: data_o = 32'h009105a3 /* 0x03cc */;
            244: data_o = 32'h00174483 /* 0x03d0 */;
            245: data_o = 32'h00910523 /* 0x03d4 */;
            246: data_o = 32'h00274483 /* 0x03d8 */;
            247: data_o = 32'h009104a3 /* 0x03dc */;
            248: data_o = 32'h00374483 /* 0x03e0 */;
            249: data_o = 32'h00910423 /* 0x03e4 */;
            250: data_o = 32'h2f8544a2 /* 0x03e8 */;
            251: data_o = 32'h24230711 /* 0x03ec */;
            252: data_o = 32'hbf81029e /* 0x03f0 */;
            253: data_o = 32'h00039563 /* 0x03f4 */;
            254: data_o = 32'hc4264304 /* 0x03f8 */;
            255: data_o = 32'he811b7f5 /* 0x03fc */;
            256: data_o = 32'h00075483 /* 0x0400 */;
            257: data_o = 32'h00911423 /* 0x0404 */;
            258: data_o = 32'h00275483 /* 0x0408 */;
            259: data_o = 32'h00911523 /* 0x040c */;
            260: data_o = 32'h4483bfe1 /* 0x0410 */;
            261: data_o = 32'h04230007 /* 0x0414 */;
            262: data_o = 32'h44830091 /* 0x0418 */;
            263: data_o = 32'h04a30017 /* 0x041c */;
            264: data_o = 32'h44830091 /* 0x0420 */;
            265: data_o = 32'h05230027 /* 0x0424 */;
            266: data_o = 32'h44830091 /* 0x0428 */;
            267: data_o = 32'h05a30037 /* 0x042c */;
            268: data_o = 32'hbf5d0091 /* 0x0430 */;
            269: data_o = 32'h01f10423 /* 0x0434 */;
            270: data_o = 32'h46014f85 /* 0x0438 */;
            271: data_o = 32'h00efd463 /* 0x043c */;
            272: data_o = 32'h0017c603 /* 0x0440 */;
            273: data_o = 32'h00c104a3 /* 0x0444 */;
            274: data_o = 32'h46014f8d /* 0x0448 */;
            275: data_o = 32'h01f71463 /* 0x044c */;
            276: data_o = 32'h0027c603 /* 0x0450 */;
            277: data_o = 32'h00c10523 /* 0x0454 */;
            278: data_o = 32'h000105a3 /* 0x0458 */;
            279: data_o = 32'h872ab72d /* 0x045c */;
            280: data_o = 32'haa95853a /* 0x0460 */;
            281: data_o = 32'h0036f713 /* 0x0464 */;
            282: data_o = 32'hc29ce319 /* 0x0468 */;
            283: data_o = 32'hf613aa4d /* 0x046c */;
            284: data_o = 32'hd71b0016 /* 0x0470 */;
            285: data_o = 32'he6110107 /* 0x0474 */;
            286: data_o = 32'h00f69023 /* 0x0478 */;
            287: data_o = 32'h00e69123 /* 0x047c */;
            288: data_o = 32'hd61baa79 /* 0x0480 */;
            289: data_o = 32'h80230087 /* 0x0484 */;
            290: data_o = 32'hd79b00f6 /* 0x0488 */;
            291: data_o = 32'h80a30187 /* 0x048c */;
            292: data_o = 32'h812300c6 /* 0x0490 */;
            293: data_o = 32'h81a300e6 /* 0x0494 */;
            294: data_o = 32'ha25100f6 /* 0x0498 */;
            295: data_o = 32'h0015071b /* 0x049c */;
            296: data_o = 32'hd61bea05 /* 0x04a0 */;
            297: data_o = 32'h80230187 /* 0x04a4 */;
            298: data_o = 32'h8be300c6 /* 0x04a8 */;
            299: data_o = 32'hd71bfae5 /* 0x04ac */;
            300: data_o = 32'h80a30107 /* 0x04b0 */;
            301: data_o = 32'h071b00e6 /* 0x04b4 */;
            302: data_o = 32'h863b0025 /* 0x04b8 */;
            303: data_o = 32'hd79b40e5 /* 0x04bc */;
            304: data_o = 32'h1fe30087 /* 0x04c0 */;
            305: data_o = 32'h8123f9c6 /* 0x04c4 */;
            306: data_o = 32'h071b00f6 /* 0x04c8 */;
            307: data_o = 32'hbf490035 /* 0x04cc */;
            308: data_o = 32'h00f68023 /* 0x04d0 */;
            309: data_o = 32'hf8e586e3 /* 0x04d4 */;
            310: data_o = 32'h0087d71b /* 0x04d8 */;
            311: data_o = 32'h00e680a3 /* 0x04dc */;
            312: data_o = 32'h0025071b /* 0x04e0 */;
            313: data_o = 32'h40e5863b /* 0x04e4 */;
            314: data_o = 32'hf7c61ce3 /* 0x04e8 */;
            315: data_o = 32'h0107d79b /* 0x04ec */;
            316: data_o = 32'hd61bbfd9 /* 0x04f0 */;
            317: data_o = 32'h80230187 /* 0x04f4 */;
            318: data_o = 32'h876300c6 /* 0x04f8 */;
            319: data_o = 32'hd71b02e5 /* 0x04fc */;
            320: data_o = 32'h80a30107 /* 0x0500 */;
            321: data_o = 32'h071b00e6 /* 0x0504 */;
            322: data_o = 32'h88630025 /* 0x0508 */;
            323: data_o = 32'hd71b00e5 /* 0x050c */;
            324: data_o = 32'h81230087 /* 0x0510 */;
            325: data_o = 32'h071b00e6 /* 0x0514 */;
            326: data_o = 32'h073b0035 /* 0x0518 */;
            327: data_o = 32'h460540e3 /* 0x051c */;
            328: data_o = 32'h00c71463 /* 0x0520 */;
            329: data_o = 32'h00f681a3 /* 0x0524 */;
            330: data_o = 32'hda088de3 /* 0x0528 */;
            331: data_o = 32'h01082783 /* 0x052c */;
            332: data_o = 32'h00083703 /* 0x0530 */;
            333: data_o = 32'h00082a23 /* 0x0534 */;
            334: data_o = 32'h8b852785 /* 0x0538 */;
            335: data_o = 32'hb355d31c /* 0x053c */;
            336: data_o = 32'h014e2783 /* 0x0540 */;
            337: data_o = 32'h27818ff9 /* 0x0544 */;
            338: data_o = 32'hbff9ffe5 /* 0x0548 */;
            339: data_o = 32'h4603571c /* 0x054c */;
            340: data_o = 32'h071b0188 /* 0x0550 */;
            341: data_o = 32'h27810015 /* 0x0554 */;
            342: data_o = 32'h8023de49 /* 0x0558 */;
            343: data_o = 32'h85e300f6 /* 0x055c */;
            344: data_o = 32'hd71bfce5 /* 0x0560 */;
            345: data_o = 32'h80a30087 /* 0x0564 */;
            346: data_o = 32'h071b00e6 /* 0x0568 */;
            347: data_o = 32'h88630025 /* 0x056c */;
            348: data_o = 32'hd71b00e5 /* 0x0570 */;
            349: data_o = 32'h81230107 /* 0x0574 */;
            350: data_o = 32'h071b00e6 /* 0x0578 */;
            351: data_o = 32'h073b0035 /* 0x057c */;
            352: data_o = 32'h460540e3 /* 0x0580 */;
            353: data_o = 32'hfac712e3 /* 0x0584 */;
            354: data_o = 32'h0187d79b /* 0x0588 */;
            355: data_o = 32'h77b3bf61 /* 0x058c */;
            356: data_o = 32'h278101d6 /* 0x0590 */;
            357: data_o = 32'hec0795e3 /* 0x0594 */;
            358: data_o = 32'hf8b578e3 /* 0x0598 */;
            359: data_o = 32'h87936789 /* 0x059c */;
            360: data_o = 32'h4b507107 /* 0x05a0 */;
            361: data_o = 32'h0086561b /* 0x05a4 */;
            362: data_o = 32'h0ff67613 /* 0x05a8 */;
            363: data_o = 32'h37fdf245 /* 0x05ac */;
            364: data_o = 32'hb511fbed /* 0x05b0 */;
            365: data_o = 32'h02fe2223 /* 0x05b4 */;
            366: data_o = 32'h01482783 /* 0x05b8 */;
            367: data_o = 32'h85e3d7b5 /* 0x05bc */;
            368: data_o = 32'hfe93f60e /* 0x05c0 */;
            369: data_o = 32'h0737001e /* 0x05c4 */;
            370: data_o = 32'h8be34000 /* 0x05c8 */;
            371: data_o = 32'h0eb7f60e /* 0x05cc */;
            372: data_o = 32'h4f0d4000 /* 0x05d0 */;
            373: data_o = 32'h37034e05 /* 0x05d4 */;
            374: data_o = 32'h4b5c0008 /* 0x05d8 */;
            375: data_o = 32'h0007861b /* 0x05dc */;
            376: data_o = 32'h0087d79b /* 0x05e0 */;
            377: data_o = 32'h0ff7f793 /* 0x05e4 */;
            378: data_o = 32'h571cd3dd /* 0x05e8 */;
            379: data_o = 32'he6b579e3 /* 0x05ec */;
            380: data_o = 32'h40a5873b /* 0x05f0 */;
            381: data_o = 32'h01884603 /* 0x05f4 */;
            382: data_o = 32'h71e32781 /* 0x05f8 */;
            383: data_o = 32'h13e3eaef /* 0x05fc */;
            384: data_o = 32'hd71be606 /* 0x0600 */;
            385: data_o = 32'h81a30087 /* 0x0604 */;
            386: data_o = 32'h812300f6 /* 0x0608 */;
            387: data_o = 32'hd71b00e6 /* 0x060c */;
            388: data_o = 32'hd79b0107 /* 0x0610 */;
            389: data_o = 32'h80a30187 /* 0x0614 */;
            390: data_o = 32'h802300e6 /* 0x0618 */;
            391: data_o = 32'h069100f6 /* 0x061c */;
            392: data_o = 32'h0045071b /* 0x0620 */;
            393: data_o = 32'h711dbd35 /* 0x0624 */;
            394: data_o = 32'h6405e8a2 /* 0x0628 */;
            395: data_o = 32'he4a6ec86 /* 0x062c */;
            396: data_o = 32'hfc4ee0ca /* 0x0630 */;
            397: data_o = 32'hf456f852 /* 0x0634 */;
            398: data_o = 32'hec5ef05a /* 0x0638 */;
            399: data_o = 32'he466e862 /* 0x063c */;
            400: data_o = 32'h0413e06a /* 0x0640 */;
            401: data_o = 32'h60638004 /* 0x0644 */;
            402: data_o = 32'h644602b4 /* 0x0648 */;
            403: data_o = 32'h64a660e6 /* 0x064c */;
            404: data_o = 32'h79e26906 /* 0x0650 */;
            405: data_o = 32'h7aa27a42 /* 0x0654 */;
            406: data_o = 32'h6be27b02 /* 0x0658 */;
            407: data_o = 32'h6ca26c42 /* 0x065c */;
            408: data_o = 32'h61256d02 /* 0x0660 */;
            409: data_o = 32'h891bb135 /* 0x0664 */;
            410: data_o = 32'h591b7ff5 /* 0x0668 */;
            411: data_o = 32'h8baa00b9 /* 0x066c */;
            412: data_o = 32'h8ab28a2e /* 0x0670 */;
            413: data_o = 32'h7c138b36 /* 0x0674 */;
            414: data_o = 32'h79930017 /* 0x0678 */;
            415: data_o = 32'h44810027 /* 0x067c */;
            416: data_o = 32'hfff90c9b /* 0x0680 */;
            417: data_o = 32'h881b8d22 /* 0x0684 */;
            418: data_o = 32'h64630004 /* 0x0688 */;
            419: data_o = 32'h45010128 /* 0x068c */;
            420: data_o = 32'h8762a0a9 /* 0x0690 */;
            421: data_o = 32'h00080663 /* 0x0694 */;
            422: data_o = 32'h93634701 /* 0x0698 */;
            423: data_o = 32'h874e010c /* 0x069c */;
            424: data_o = 32'h80000793 /* 0x06a0 */;
            425: data_o = 32'h030787bb /* 0x06a4 */;
            426: data_o = 32'h014786bb /* 0x06a8 */;
            427: data_o = 32'h736387b6 /* 0x06ac */;
            428: data_o = 32'h87ea00d4 /* 0x06b0 */;
            429: data_o = 32'h0007859b /* 0x06b4 */;
            430: data_o = 32'h85634601 /* 0x06b8 */;
            431: data_o = 32'h9613000a /* 0x06bc */;
            432: data_o = 32'h96560084 /* 0x06c0 */;
            433: data_o = 32'h05634681 /* 0x06c4 */;
            434: data_o = 32'h9693000b /* 0x06c8 */;
            435: data_o = 32'h96da0084 /* 0x06cc */;
            436: data_o = 32'hf0ef855e /* 0x06d0 */;
            437: data_o = 32'h0485bbff /* 0x06d4 */;
            438: data_o = 32'h60e6d55d /* 0x06d8 */;
            439: data_o = 32'h64a66446 /* 0x06dc */;
            440: data_o = 32'h79e26906 /* 0x06e0 */;
            441: data_o = 32'h7aa27a42 /* 0x06e4 */;
            442: data_o = 32'h6be27b02 /* 0x06e8 */;
            443: data_o = 32'h6ca26c42 /* 0x06ec */;
            444: data_o = 32'h61256d02 /* 0x06f0 */;
            445: data_o = 32'h71798082 /* 0x06f4 */;
            446: data_o = 32'hf022f406 /* 0x06f8 */;
            447: data_o = 32'he84aec26 /* 0x06fc */;
            448: data_o = 32'h00010623 /* 0x0700 */;
            449: data_o = 32'hceb14781 /* 0x0704 */;
            450: data_o = 32'h00800737 /* 0x0708 */;
            451: data_o = 32'hfa6357fd /* 0x070c */;
            452: data_o = 32'h073704e5 /* 0x0710 */;
            453: data_o = 32'h84360010 /* 0x0714 */;
            454: data_o = 32'h04e6f563 /* 0x0718 */;
            455: data_o = 32'h0095959b /* 0x071c */;
            456: data_o = 32'h042347cd /* 0x0720 */;
            457: data_o = 32'hd79b00f1 /* 0x0724 */;
            458: data_o = 32'h04a30185 /* 0x0728 */;
            459: data_o = 32'hd79b00f1 /* 0x072c */;
            460: data_o = 32'hd59b0105 /* 0x0730 */;
            461: data_o = 32'h89320085 /* 0x0734 */;
            462: data_o = 32'h00b105a3 /* 0x0738 */;
            463: data_o = 32'h46814705 /* 0x073c */;
            464: data_o = 32'h05930030 /* 0x0740 */;
            465: data_o = 32'h05230280 /* 0x0744 */;
            466: data_o = 32'h84aa00f1 /* 0x0748 */;
            467: data_o = 32'hedbff0ef /* 0x074c */;
            468: data_o = 32'h00c4159b /* 0x0750 */;
            469: data_o = 32'h86ca4709 /* 0x0754 */;
            470: data_o = 32'h85264601 /* 0x0758 */;
            471: data_o = 32'hecbff0ef /* 0x075c */;
            472: data_o = 32'h70a287aa /* 0x0760 */;
            473: data_o = 32'h64e27402 /* 0x0764 */;
            474: data_o = 32'h853e6942 /* 0x0768 */;
            475: data_o = 32'h80826145 /* 0x076c */;
            476: data_o = 32'h4785b759 /* 0x0770 */;
            477: data_o = 32'h00b797bb /* 0x0774 */;
            478: data_o = 32'hfff7c793 /* 0x0778 */;
            479: data_o = 32'h163b8fe9 /* 0x077c */;
            480: data_o = 32'h8fd100b6 /* 0x0780 */;
            481: data_o = 32'h0007851b /* 0x0784 */;
            482: data_o = 32'h71798082 /* 0x0788 */;
            483: data_o = 32'hf406e84a /* 0x078c */;
            484: data_o = 32'hec26f022 /* 0x0790 */;
            485: data_o = 32'h892ae44e /* 0x0794 */;
            486: data_o = 32'hcd254789 /* 0x0798 */;
            487: data_o = 32'h8436852e /* 0x079c */;
            488: data_o = 32'h071bc699 /* 0x07a0 */;
            489: data_o = 32'h4689ffd6 /* 0x07a4 */;
            490: data_o = 32'hf4634789 /* 0x07a8 */;
            491: data_o = 32'h478906e6 /* 0x07ac */;
            492: data_o = 32'h02f60263 /* 0x07b0 */;
            493: data_o = 32'h0663478d /* 0x07b4 */;
            494: data_o = 32'h079306f6 /* 0x07b8 */;
            495: data_o = 32'h3633fff6 /* 0x07bc */;
            496: data_o = 32'h448100f0 /* 0x07c0 */;
            497: data_o = 32'heb914981 /* 0x07c4 */;
            498: data_o = 32'h0004071b /* 0x07c8 */;
            499: data_o = 32'h4789c499 /* 0x07cc */;
            500: data_o = 32'ha081c709 /* 0x07d0 */;
            501: data_o = 32'h49854481 /* 0x07d4 */;
            502: data_o = 32'h45a14601 /* 0x07d8 */;
            503: data_o = 32'hf97ff0ef /* 0x07dc */;
            504: data_o = 32'h45a5864e /* 0x07e0 */;
            505: data_o = 32'hf0ef2501 /* 0x07e4 */;
            506: data_o = 32'h8626f8df /* 0x07e8 */;
            507: data_o = 32'h250145a9 /* 0x07ec */;
            508: data_o = 32'hf83ff0ef /* 0x07f0 */;
            509: data_o = 32'h45ad4601 /* 0x07f4 */;
            510: data_o = 32'hf0ef2501 /* 0x07f8 */;
            511: data_o = 32'h8622f79f /* 0x07fc */;
            512: data_o = 32'h250145b1 /* 0x0800 */;
            513: data_o = 32'hf6fff0ef /* 0x0804 */;
            514: data_o = 32'h00093783 /* 0x0808 */;
            515: data_o = 32'hcfc82501 /* 0x080c */;
            516: data_o = 32'h70a24781 /* 0x0810 */;
            517: data_o = 32'h64e27402 /* 0x0814 */;
            518: data_o = 32'h69a26942 /* 0x0818 */;
            519: data_o = 32'h6145853e /* 0x081c */;
            520: data_o = 32'h44858082 /* 0x0820 */;
            521: data_o = 32'h46014981 /* 0x0824 */;
            522: data_o = 32'h8163b745 /* 0x0828 */;
            523: data_o = 32'h711d1c06 /* 0x082c */;
            524: data_o = 32'hec86e8a2 /* 0x0830 */;
            525: data_o = 32'he0cae4a6 /* 0x0834 */;
            526: data_o = 32'hf852fc4e /* 0x0838 */;
            527: data_o = 32'hf05af456 /* 0x083c */;
            528: data_o = 32'he862ec5e /* 0x0840 */;
            529: data_o = 32'he06ae466 /* 0x0844 */;
            530: data_o = 32'h00b6e7b3 /* 0x0848 */;
            531: data_o = 32'h0ff00713 /* 0x084c */;
            532: data_o = 32'h557d842a /* 0x0850 */;
            533: data_o = 32'h16f76663 /* 0x0854 */;
            534: data_o = 32'h949b8b32 /* 0x0858 */;
            535: data_o = 32'h999b0095 /* 0x085c */;
            536: data_o = 32'h4a810036 /* 0x0860 */;
            537: data_o = 32'h6c414a01 /* 0x0864 */;
            538: data_o = 32'h03f00c93 /* 0x0868 */;
            539: data_o = 32'h09134d21 /* 0x086c */;
            540: data_o = 32'he4630a00 /* 0x0870 */;
            541: data_o = 32'h09130184 /* 0x0874 */;
            542: data_o = 32'h46850a80 /* 0x0878 */;
            543: data_o = 32'h85ca4601 /* 0x087c */;
            544: data_o = 32'hf0ef8522 /* 0x0880 */;
            545: data_o = 32'h2501f09f /* 0x0884 */;
            546: data_o = 32'h5575c501 /* 0x0888 */;
            547: data_o = 32'h917ff06f /* 0x088c */;
            548: data_o = 32'h0084d59b /* 0x0890 */;
            549: data_o = 32'h46054685 /* 0x0894 */;
            550: data_o = 32'h0ff5f593 /* 0x0898 */;
            551: data_o = 32'hf0ef8522 /* 0x089c */;
            552: data_o = 32'h2501eedf /* 0x08a0 */;
            553: data_o = 32'h5575c501 /* 0x08a4 */;
            554: data_o = 32'h8fbff06f /* 0x08a8 */;
            555: data_o = 32'h46094685 /* 0x08ac */;
            556: data_o = 32'h0ff4f593 /* 0x08b0 */;
            557: data_o = 32'hf0ef8522 /* 0x08b4 */;
            558: data_o = 32'h2501ed5f /* 0x08b8 */;
            559: data_o = 32'h5575c501 /* 0x08bc */;
            560: data_o = 32'h8e3ff06f /* 0x08c0 */;
            561: data_o = 32'h46014685 /* 0x08c4 */;
            562: data_o = 32'h00196593 /* 0x08c8 */;
            563: data_o = 32'hf0ef8522 /* 0x08cc */;
            564: data_o = 32'h2501ebdf /* 0x08d0 */;
            565: data_o = 32'h5575c501 /* 0x08d4 */;
            566: data_o = 32'h8cbff06f /* 0x08d8 */;
            567: data_o = 32'h460d4681 /* 0x08dc */;
            568: data_o = 32'h04000593 /* 0x08e0 */;
            569: data_o = 32'hf0ef8522 /* 0x08e4 */;
            570: data_o = 32'h2501ea5f /* 0x08e8 */;
            571: data_o = 32'h5575c501 /* 0x08ec */;
            572: data_o = 32'h8b3ff06f /* 0x08f0 */;
            573: data_o = 32'h0e041463 /* 0x08f4 */;
            574: data_o = 32'hf06f5575 /* 0x08f8 */;
            575: data_o = 32'hfbe38a9f /* 0x08fc */;
            576: data_o = 32'h9913ff4c /* 0x0900 */;
            577: data_o = 32'h995a006a /* 0x0904 */;
            578: data_o = 32'h85ca4b81 /* 0x0908 */;
            579: data_o = 32'hf0ef8522 /* 0x090c */;
            580: data_o = 32'h25018bdf /* 0x0910 */;
            581: data_o = 32'h5575c501 /* 0x0914 */;
            582: data_o = 32'h88bff06f /* 0x0918 */;
            583: data_o = 32'h00190593 /* 0x091c */;
            584: data_o = 32'hf0ef8522 /* 0x0920 */;
            585: data_o = 32'h25018a9f /* 0x0924 */;
            586: data_o = 32'h5575c501 /* 0x0928 */;
            587: data_o = 32'h877ff06f /* 0x092c */;
            588: data_o = 32'h00290593 /* 0x0930 */;
            589: data_o = 32'hf0ef8522 /* 0x0934 */;
            590: data_o = 32'h2501895f /* 0x0938 */;
            591: data_o = 32'h5575c501 /* 0x093c */;
            592: data_o = 32'h863ff06f /* 0x0940 */;
            593: data_o = 32'h00390593 /* 0x0944 */;
            594: data_o = 32'hf0ef8522 /* 0x0948 */;
            595: data_o = 32'h2501881f /* 0x094c */;
            596: data_o = 32'h5575c501 /* 0x0950 */;
            597: data_o = 32'h84fff06f /* 0x0954 */;
            598: data_o = 32'h00490593 /* 0x0958 */;
            599: data_o = 32'hf0ef8522 /* 0x095c */;
            600: data_o = 32'h250186df /* 0x0960 */;
            601: data_o = 32'h5575c501 /* 0x0964 */;
            602: data_o = 32'h83bff06f /* 0x0968 */;
            603: data_o = 32'h00590593 /* 0x096c */;
            604: data_o = 32'hf0ef8522 /* 0x0970 */;
            605: data_o = 32'h2501859f /* 0x0974 */;
            606: data_o = 32'h5575c501 /* 0x0978 */;
            607: data_o = 32'h827ff06f /* 0x097c */;
            608: data_o = 32'h00690593 /* 0x0980 */;
            609: data_o = 32'hf0ef8522 /* 0x0984 */;
            610: data_o = 32'h2501845f /* 0x0988 */;
            611: data_o = 32'h5575c501 /* 0x098c */;
            612: data_o = 32'h813ff06f /* 0x0990 */;
            613: data_o = 32'h00790593 /* 0x0994 */;
            614: data_o = 32'hf0ef8522 /* 0x0998 */;
            615: data_o = 32'h2501831f /* 0x099c */;
            616: data_o = 32'h5575c501 /* 0x09a0 */;
            617: data_o = 32'hffeff06f /* 0x09a4 */;
            618: data_o = 32'h09212b85 /* 0x09a8 */;
            619: data_o = 32'hf5ab9fe3 /* 0x09ac */;
            620: data_o = 32'h879b0a85 /* 0x09b0 */;
            621: data_o = 32'h849b000a /* 0x09b4 */;
            622: data_o = 32'heae30404 /* 0x09b8 */;
            623: data_o = 32'h4501eb37 /* 0x09bc */;
            624: data_o = 32'h644660e6 /* 0x09c0 */;
            625: data_o = 32'h690664a6 /* 0x09c4 */;
            626: data_o = 32'h7a4279e2 /* 0x09c8 */;
            627: data_o = 32'h7b027aa2 /* 0x09cc */;
            628: data_o = 32'h6c426be2 /* 0x09d0 */;
            629: data_o = 32'h6d026ca2 /* 0x09d4 */;
            630: data_o = 32'h80826125 /* 0x09d8 */;
            631: data_o = 32'haa03601c /* 0x09dc */;
            632: data_o = 32'h5a1b0247 /* 0x09e0 */;
            633: data_o = 32'h7a13010a /* 0x09e4 */;
            634: data_o = 32'hbf1107fa /* 0x09e8 */;
            635: data_o = 32'h80824501 /* 0x09ec */;
            636: data_o = 32'h711dbd2d /* 0x09f0 */;
            637: data_o = 32'he0cae4a6 /* 0x09f4 */;
            638: data_o = 32'hf852fc4e /* 0x09f8 */;
            639: data_o = 32'hf05af456 /* 0x09fc */;
            640: data_o = 32'h89beec5e /* 0x0a00 */;
            641: data_o = 32'he8a2ec86 /* 0x0a04 */;
            642: data_o = 32'he466e862 /* 0x0a08 */;
            643: data_o = 32'h00387793 /* 0x0a0c */;
            644: data_o = 32'h8b2e8aaa /* 0x0a10 */;
            645: data_o = 32'h8bb68932 /* 0x0a14 */;
            646: data_o = 32'h8a4284ba /* 0x0a18 */;
            647: data_o = 32'h8432c3b5 /* 0x0a1c */;
            648: data_o = 32'h85229426 /* 0x0a20 */;
            649: data_o = 32'h40940633 /* 0x0a24 */;
            650: data_o = 32'h7a13e4a5 /* 0x0a28 */;
            651: data_o = 32'h0b63002a /* 0x0a2c */;
            652: data_o = 32'h1982000a /* 0x0a30 */;
            653: data_o = 32'h41240433 /* 0x0a34 */;
            654: data_o = 32'h0209d993 /* 0x0a38 */;
            655: data_o = 32'h00890533 /* 0x0a3c */;
            656: data_o = 32'h07346163 /* 0x0a40 */;
            657: data_o = 32'h644660e6 /* 0x0a44 */;
            658: data_o = 32'h690664a6 /* 0x0a48 */;
            659: data_o = 32'h7a4279e2 /* 0x0a4c */;
            660: data_o = 32'h7b027aa2 /* 0x0a50 */;
            661: data_o = 32'h6c426be2 /* 0x0a54 */;
            662: data_o = 32'h61256ca2 /* 0x0a58 */;
            663: data_o = 32'h56fd8082 /* 0x0a5c */;
            664: data_o = 32'h051385da /* 0x0a60 */;
            665: data_o = 32'h9a820200 /* 0x0a64 */;
            666: data_o = 32'h86330405 /* 0x0a68 */;
            667: data_o = 32'h68e3008c /* 0x0a6c */;
            668: data_o = 32'h4401ff84 /* 0x0a70 */;
            669: data_o = 32'h009c6463 /* 0x0a74 */;
            670: data_o = 32'h409c0433 /* 0x0a78 */;
            671: data_o = 32'hb74d944a /* 0x0a7c */;
            672: data_o = 32'h02099c13 /* 0x0a80 */;
            673: data_o = 32'h0cb3843a /* 0x0a84 */;
            674: data_o = 32'h5c1340e6 /* 0x0a88 */;
            675: data_o = 32'hbff1020c /* 0x0a8c */;
            676: data_o = 32'h87b314fd /* 0x0a90 */;
            677: data_o = 32'hc503009b /* 0x0a94 */;
            678: data_o = 32'h56fd0007 /* 0x0a98 */;
            679: data_o = 32'h9a8285da /* 0x0a9c */;
            680: data_o = 32'h862ab749 /* 0x0aa0 */;
            681: data_o = 32'h85da56fd /* 0x0aa4 */;
            682: data_o = 32'h02000513 /* 0x0aa8 */;
            683: data_o = 32'h04059a82 /* 0x0aac */;
            684: data_o = 32'h7179b771 /* 0x0ab0 */;
            685: data_o = 32'hf022f406 /* 0x0ab4 */;
            686: data_o = 32'h8ec28e3e /* 0x0ab8 */;
            687: data_o = 32'h584287c6 /* 0x0abc */;
            688: data_o = 32'h7813e299 /* 0x0ac0 */;
            689: data_o = 32'h7293fef8 /* 0x0ac4 */;
            690: data_o = 32'h83634008 /* 0x0ac8 */;
            691: data_o = 32'hc6a10002 /* 0x0acc */;
            692: data_o = 32'h02087313 /* 0x0ad0 */;
            693: data_o = 32'h06100893 /* 0x0ad4 */;
            694: data_o = 32'h00030463 /* 0x0ad8 */;
            695: data_o = 32'h04100893 /* 0x0adc */;
            696: data_o = 32'h8f8a8f36 /* 0x0ae0 */;
            697: data_o = 32'h44254681 /* 0x0ae4 */;
            698: data_o = 32'h009338d9 /* 0x0ae8 */;
            699: data_o = 32'h73b30200 /* 0x0aec */;
            700: data_o = 32'hf31303cf /* 0x0af0 */;
            701: data_o = 32'h6b630ff3 /* 0x0af4 */;
            702: data_o = 32'h031b0474 /* 0x0af8 */;
            703: data_o = 32'h73130303 /* 0x0afc */;
            704: data_o = 32'h80230ff3 /* 0x0b00 */;
            705: data_o = 32'h0685006f /* 0x0b04 */;
            706: data_o = 32'h03cf5333 /* 0x0b08 */;
            707: data_o = 32'h01cf6563 /* 0x0b0c */;
            708: data_o = 32'h9b630f85 /* 0x0b10 */;
            709: data_o = 32'h73130216 /* 0x0b14 */;
            710: data_o = 32'h88c20028 /* 0x0b18 */;
            711: data_o = 32'h06031163 /* 0x0b1c */;
            712: data_o = 32'h00187313 /* 0x0b20 */;
            713: data_o = 32'h0863cb89 /* 0x0b24 */;
            714: data_o = 32'he7090003 /* 0x0b28 */;
            715: data_o = 32'h00c8f893 /* 0x0b2c */;
            716: data_o = 32'h00088363 /* 0x0b30 */;
            717: data_o = 32'h9f1337fd /* 0x0b34 */;
            718: data_o = 32'h5f13020e /* 0x0b38 */;
            719: data_o = 32'h0893020f /* 0x0b3c */;
            720: data_o = 32'h0f930200 /* 0x0b40 */;
            721: data_o = 32'ha8190300 /* 0x0b44 */;
            722: data_o = 32'hb7558f1a /* 0x0b48 */;
            723: data_o = 32'h0068833b /* 0x0b4c */;
            724: data_o = 32'h03b3b77d /* 0x0b50 */;
            725: data_o = 32'h802300d1 /* 0x0b54 */;
            726: data_o = 32'h068501f3 /* 0x0b58 */;
            727: data_o = 32'h01e6f463 /* 0x0b5c */;
            728: data_o = 32'hff1699e3 /* 0x0b60 */;
            729: data_o = 32'h02079f13 /* 0x0b64 */;
            730: data_o = 32'h020f5f13 /* 0x0b68 */;
            731: data_o = 32'h0f9348fd /* 0x0b6c */;
            732: data_o = 32'h06630300 /* 0x0b70 */;
            733: data_o = 32'hf4630003 /* 0x0b74 */;
            734: data_o = 32'hfa6301e6 /* 0x0b78 */;
            735: data_o = 32'h789304d8 /* 0x0b7c */;
            736: data_o = 32'h8c630108 /* 0x0b80 */;
            737: data_o = 32'h9b630808 /* 0x0b84 */;
            738: data_o = 32'hcaa90402 /* 0x0b88 */;
            739: data_o = 32'hde931e82 /* 0x0b8c */;
            740: data_o = 32'h8863020e /* 0x0b90 */;
            741: data_o = 32'h989301d6 /* 0x0b94 */;
            742: data_o = 32'hd8930207 /* 0x0b98 */;
            743: data_o = 32'h9f630208 /* 0x0b9c */;
            744: data_o = 32'h88930316 /* 0x0ba0 */;
            745: data_o = 32'h8a63fff6 /* 0x0ba4 */;
            746: data_o = 32'h43410208 /* 0x0ba8 */;
            747: data_o = 32'h0a6316f9 /* 0x0bac */;
            748: data_o = 32'h86c6026e /* 0x0bb0 */;
            749: data_o = 32'h16634889 /* 0x0bb4 */;
            750: data_o = 32'h48fd051e /* 0x0bb8 */;
            751: data_o = 32'h06d8eb63 /* 0x0bbc */;
            752: data_o = 32'h02068413 /* 0x0bc0 */;
            753: data_o = 32'h002408b3 /* 0x0bc4 */;
            754: data_o = 32'h06200313 /* 0x0bc8 */;
            755: data_o = 32'h03b3a805 /* 0x0bcc */;
            756: data_o = 32'h802300d1 /* 0x0bd0 */;
            757: data_o = 32'h068501f3 /* 0x0bd4 */;
            758: data_o = 32'h4681bf69 /* 0x0bd8 */;
            759: data_o = 32'h1be348c1 /* 0x0bdc */;
            760: data_o = 32'h7893fd1e /* 0x0be0 */;
            761: data_o = 32'h9e630208 /* 0x0be4 */;
            762: data_o = 32'h48fd0408 /* 0x0be8 */;
            763: data_o = 32'h04d8e363 /* 0x0bec */;
            764: data_o = 32'h02068413 /* 0x0bf0 */;
            765: data_o = 32'h002408b3 /* 0x0bf4 */;
            766: data_o = 32'h07800313 /* 0x0bf8 */;
            767: data_o = 32'hfe688023 /* 0x0bfc */;
            768: data_o = 32'h48fd0685 /* 0x0c00 */;
            769: data_o = 32'h02d8e763 /* 0x0c04 */;
            770: data_o = 32'h02068413 /* 0x0c08 */;
            771: data_o = 32'h002408b3 /* 0x0c0c */;
            772: data_o = 32'h03000313 /* 0x0c10 */;
            773: data_o = 32'hfe688023 /* 0x0c14 */;
            774: data_o = 32'h48fd0685 /* 0x0c18 */;
            775: data_o = 32'h00d8eb63 /* 0x0c1c */;
            776: data_o = 32'h8713cb1d /* 0x0c20 */;
            777: data_o = 32'h970a0206 /* 0x0c24 */;
            778: data_o = 32'h02d00893 /* 0x0c28 */;
            779: data_o = 32'hff170023 /* 0x0c2c */;
            780: data_o = 32'h87360685 /* 0x0c30 */;
            781: data_o = 32'hf0ef868a /* 0x0c34 */;
            782: data_o = 32'h70a2dbdf /* 0x0c38 */;
            783: data_o = 32'h61457402 /* 0x0c3c */;
            784: data_o = 32'h48fd8082 /* 0x0c40 */;
            785: data_o = 32'hfed8e7e3 /* 0x0c44 */;
            786: data_o = 32'h02068413 /* 0x0c48 */;
            787: data_o = 32'h002408b3 /* 0x0c4c */;
            788: data_o = 32'h05800313 /* 0x0c50 */;
            789: data_o = 32'h7713b765 /* 0x0c54 */;
            790: data_o = 32'hc7190048 /* 0x0c58 */;
            791: data_o = 32'h02068713 /* 0x0c5c */;
            792: data_o = 32'h0893970a /* 0x0c60 */;
            793: data_o = 32'hb7d902b0 /* 0x0c64 */;
            794: data_o = 32'h00887713 /* 0x0c68 */;
            795: data_o = 32'h8713d379 /* 0x0c6c */;
            796: data_o = 32'h970a0206 /* 0x0c70 */;
            797: data_o = 32'h02000893 /* 0x0c74 */;
            798: data_o = 32'h711dbf55 /* 0x0c78 */;
            799: data_o = 32'h84bee4a6 /* 0x0c7c */;
            800: data_o = 32'ha2a527d3 /* 0x0c80 */;
            801: data_o = 32'hfc4ee0ca /* 0x0c84 */;
            802: data_o = 32'hf05af852 /* 0x0c88 */;
            803: data_o = 32'he8a2ec86 /* 0x0c8c */;
            804: data_o = 32'hec5ef456 /* 0x0c90 */;
            805: data_o = 32'h8a2e892a /* 0x0c94 */;
            806: data_o = 32'h8b3a89b2 /* 0x0c98 */;
            807: data_o = 32'h1797cf99 /* 0x0c9c */;
            808: data_o = 32'hb7870000 /* 0x0ca0 */;
            809: data_o = 32'h97d37f27 /* 0x0ca4 */;
            810: data_o = 32'heb81a2a7 /* 0x0ca8 */;
            811: data_o = 32'h00001797 /* 0x0cac */;
            812: data_o = 32'h7ec7b787 /* 0x0cb0 */;
            813: data_o = 32'ha2f517d3 /* 0x0cb4 */;
            814: data_o = 32'h6446c38d /* 0x0cb8 */;
            815: data_o = 32'h7aa260e6 /* 0x0cbc */;
            816: data_o = 32'h87a66be2 /* 0x0cc0 */;
            817: data_o = 32'h64a6875a /* 0x0cc4 */;
            818: data_o = 32'h864e7b02 /* 0x0cc8 */;
            819: data_o = 32'h79e285d2 /* 0x0ccc */;
            820: data_o = 32'h854a7a42 /* 0x0cd0 */;
            821: data_o = 32'h61256906 /* 0x0cd4 */;
            822: data_o = 32'h07d3acb1 /* 0x0cd8 */;
            823: data_o = 32'h17d3f200 /* 0x0cdc */;
            824: data_o = 32'h17d3a2f5 /* 0x0ce0 */;
            825: data_o = 32'h865322a5 /* 0x0ce4 */;
            826: data_o = 32'he399e207 /* 0x0ce8 */;
            827: data_o = 32'he2050653 /* 0x0cec */;
            828: data_o = 32'h4004f713 /* 0x0cf0 */;
            829: data_o = 32'h4699e311 /* 0x0cf4 */;
            830: data_o = 32'h03465793 /* 0x0cf8 */;
            831: data_o = 32'h7ff7f793 /* 0x0cfc */;
            832: data_o = 32'hc017879b /* 0x0d00 */;
            833: data_o = 32'hd2078753 /* 0x0d04 */;
            834: data_o = 32'h00001797 /* 0x0d08 */;
            835: data_o = 32'h7987b687 /* 0x0d0c */;
            836: data_o = 32'h00001797 /* 0x0d10 */;
            837: data_o = 32'h7987b787 /* 0x0d14 */;
            838: data_o = 32'h3ff00593 /* 0x0d18 */;
            839: data_o = 32'h00c61793 /* 0x0d1c */;
            840: data_o = 32'h83b115d2 /* 0x0d20 */;
            841: data_o = 32'h15978fcd /* 0x0d24 */;
            842: data_o = 32'h77430000 /* 0x0d28 */;
            843: data_o = 32'h86d37ad7 /* 0x0d2c */;
            844: data_o = 32'hb787f207 /* 0x0d30 */;
            845: data_o = 32'h179778a5 /* 0x0d34 */;
            846: data_o = 32'h15170000 /* 0x0d38 */;
            847: data_o = 32'hf7d30000 /* 0x0d3c */;
            848: data_o = 32'hb6870af6 /* 0x0d40 */;
            849: data_o = 32'h17977827 /* 0x0d44 */;
            850: data_o = 32'hf7c30000 /* 0x0d48 */;
            851: data_o = 32'h95d372d7 /* 0x0d4c */;
            852: data_o = 32'hb787c207 /* 0x0d50 */;
            853: data_o = 32'h179777a7 /* 0x0d54 */;
            854: data_o = 32'hb7070000 /* 0x0d58 */;
            855: data_o = 32'h86d37727 /* 0x0d5c */;
            856: data_o = 32'h8b9bd205 /* 0x0d60 */;
            857: data_o = 32'hf7c30005 /* 0x0d64 */;
            858: data_o = 32'h370772f6 /* 0x0d68 */;
            859: data_o = 32'h15177965 /* 0x0d6c */;
            860: data_o = 32'h97d30000 /* 0x0d70 */;
            861: data_o = 32'h87d3c207 /* 0x0d74 */;
            862: data_o = 32'h879bd207 /* 0x0d78 */;
            863: data_o = 32'h17d23ff7 /* 0x0d7c */;
            864: data_o = 32'h12e7f7d3 /* 0x0d80 */;
            865: data_o = 32'h76a53707 /* 0x0d84 */;
            866: data_o = 32'h00001517 /* 0x0d88 */;
            867: data_o = 32'h7ae6f6c7 /* 0x0d8c */;
            868: data_o = 32'h75853707 /* 0x0d90 */;
            869: data_o = 32'h00001517 /* 0x0d94 */;
            870: data_o = 32'h75453587 /* 0x0d98 */;
            871: data_o = 32'h00001517 /* 0x0d9c */;
            872: data_o = 32'h75453007 /* 0x0da0 */;
            873: data_o = 32'h00001517 /* 0x0da4 */;
            874: data_o = 32'h12d6f653 /* 0x0da8 */;
            875: data_o = 32'h02d6f7d3 /* 0x0dac */;
            876: data_o = 32'h1ae67753 /* 0x0db0 */;
            877: data_o = 32'h02b77753 /* 0x0db4 */;
            878: data_o = 32'h1ae67753 /* 0x0db8 */;
            879: data_o = 32'h02077753 /* 0x0dbc */;
            880: data_o = 32'h1ae67653 /* 0x0dc0 */;
            881: data_o = 32'h75453707 /* 0x0dc4 */;
            882: data_o = 32'h00001517 /* 0x0dc8 */;
            883: data_o = 32'h0ad77753 /* 0x0dcc */;
            884: data_o = 32'h02e67653 /* 0x0dd0 */;
            885: data_o = 32'h73853707 /* 0x0dd4 */;
            886: data_o = 32'h1ac7f7d3 /* 0x0dd8 */;
            887: data_o = 32'h02e7f7d3 /* 0x0ddc */;
            888: data_o = 32'hf2078753 /* 0x0de0 */;
            889: data_o = 32'h12e7f7d3 /* 0x0de4 */;
            890: data_o = 32'he20787d3 /* 0x0de8 */;
            891: data_o = 32'hf20607d3 /* 0x0dec */;
            892: data_o = 32'hf2078753 /* 0x0df0 */;
            893: data_o = 32'ha2e79553 /* 0x0df4 */;
            894: data_o = 32'h77d3c519 /* 0x0df8 */;
            895: data_o = 32'h8b9b1ab7 /* 0x0dfc */;
            896: data_o = 32'h87d3fff5 /* 0x0e00 */;
            897: data_o = 32'h0593e207 /* 0x0e04 */;
            898: data_o = 32'h841b0c60 /* 0x0e08 */;
            899: data_o = 32'hb433063b /* 0x0e0c */;
            900: data_o = 32'hd5930085 /* 0x0e10 */;
            901: data_o = 32'h898500b4 /* 0x0e14 */;
            902: data_o = 32'hcd950411 /* 0x0e18 */;
            903: data_o = 32'h00001597 /* 0x0e1c */;
            904: data_o = 32'h6ec5b787 /* 0x0e20 */;
            905: data_o = 32'hf2060753 /* 0x0e24 */;
            906: data_o = 32'ha2e785d3 /* 0x0e28 */;
            907: data_o = 32'h1597c9ed /* 0x0e2c */;
            908: data_o = 32'hb7870000 /* 0x0e30 */;
            909: data_o = 32'h15d36e25 /* 0x0e34 */;
            910: data_o = 32'hc1f5a2f7 /* 0x0e38 */;
            911: data_o = 32'h0006871b /* 0x0e3c */;
            912: data_o = 32'hd6634681 /* 0x0e40 */;
            913: data_o = 32'h073b00eb /* 0x0e44 */;
            914: data_o = 32'h069b4177 /* 0x0e48 */;
            915: data_o = 32'he493fff7 /* 0x0e4c */;
            916: data_o = 32'h44014004 /* 0x0e50 */;
            917: data_o = 32'h47014b81 /* 0x0e54 */;
            918: data_o = 32'h01647463 /* 0x0e58 */;
            919: data_o = 32'h408b073b /* 0x0e5c */;
            920: data_o = 32'h0024fa93 /* 0x0e60 */;
            921: data_o = 32'h000a8463 /* 0x0e64 */;
            922: data_o = 32'h4701c011 /* 0x0e68 */;
            923: data_o = 32'h000b8a63 /* 0x0e6c */;
            924: data_o = 32'hf20607d3 /* 0x0e70 */;
            925: data_o = 32'hf2078753 /* 0x0e74 */;
            926: data_o = 32'h1ae7f7d3 /* 0x0e78 */;
            927: data_o = 32'he2078653 /* 0x0e7c */;
            928: data_o = 32'hf20007d3 /* 0x0e80 */;
            929: data_o = 32'ha2f517d3 /* 0x0e84 */;
            930: data_o = 32'h07d3c799 /* 0x0e88 */;
            931: data_o = 32'h97d3f206 /* 0x0e8c */;
            932: data_o = 32'h865322f7 /* 0x0e90 */;
            933: data_o = 32'h0553e207 /* 0x0e94 */;
            934: data_o = 32'h77fdf206 /* 0x0e98 */;
            935: data_o = 32'h7ff78793 /* 0x0e9c */;
            936: data_o = 32'h8fe5864e /* 0x0ea0 */;
            937: data_o = 32'h854a85d2 /* 0x0ea4 */;
            938: data_o = 32'h08c000ef /* 0x0ea8 */;
            939: data_o = 32'hcc21862a /* 0x0eac */;
            940: data_o = 32'h0204f493 /* 0x0eb0 */;
            941: data_o = 32'h04500513 /* 0x0eb4 */;
            942: data_o = 32'h0513e099 /* 0x0eb8 */;
            943: data_o = 32'h56fd0650 /* 0x0ebc */;
            944: data_o = 32'h049385d2 /* 0x0ec0 */;
            945: data_o = 32'h99020016 /* 0x0ec4 */;
            946: data_o = 32'h41fbd69b /* 0x0ec8 */;
            947: data_o = 32'h00dbc633 /* 0x0ecc */;
            948: data_o = 32'he03e4795 /* 0x0ed0 */;
            949: data_o = 32'h40d606bb /* 0x0ed4 */;
            950: data_o = 32'hfff4089b /* 0x0ed8 */;
            951: data_o = 32'h48018626 /* 0x0edc */;
            952: data_o = 32'hd71b47a9 /* 0x0ee0 */;
            953: data_o = 32'h85d201fb /* 0x0ee4 */;
            954: data_o = 32'hf0ef854a /* 0x0ee8 */;
            955: data_o = 32'h862abc9f /* 0x0eec */;
            956: data_o = 32'h000a8b63 /* 0x0ef0 */;
            957: data_o = 32'h04331b02 /* 0x0ef4 */;
            958: data_o = 32'h5b134135 /* 0x0ef8 */;
            959: data_o = 32'h8633020b /* 0x0efc */;
            960: data_o = 32'h62630089 /* 0x0f00 */;
            961: data_o = 32'h60e60364 /* 0x0f04 */;
            962: data_o = 32'h64a66446 /* 0x0f08 */;
            963: data_o = 32'h79e26906 /* 0x0f0c */;
            964: data_o = 32'h7aa27a42 /* 0x0f10 */;
            965: data_o = 32'h6be27b02 /* 0x0f14 */;
            966: data_o = 32'h61258532 /* 0x0f18 */;
            967: data_o = 32'hde858082 /* 0x0f1c */;
            968: data_o = 32'h36fddb1d /* 0x0f20 */;
            969: data_o = 32'h56fdbf0d /* 0x0f24 */;
            970: data_o = 32'h051385d2 /* 0x0f28 */;
            971: data_o = 32'h99020200 /* 0x0f2c */;
            972: data_o = 32'hb7f10405 /* 0x0f30 */;
            973: data_o = 32'h27d3883e /* 0x0f34 */;
            974: data_o = 32'heb81a2a5 /* 0x0f38 */;
            975: data_o = 32'h00001697 /* 0x0f3c */;
            976: data_o = 32'h869387ba /* 0x0f40 */;
            977: data_o = 32'h470d2cc6 /* 0x0f44 */;
            978: data_o = 32'h1797b46d /* 0x0f48 */;
            979: data_o = 32'hb7870000 /* 0x0f4c */;
            980: data_o = 32'h17d354e7 /* 0x0f50 */;
            981: data_o = 32'hcb81a2f5 /* 0x0f54 */;
            982: data_o = 32'h00001697 /* 0x0f58 */;
            983: data_o = 32'h869387ba /* 0x0f5c */;
            984: data_o = 32'h47112b86 /* 0x0f60 */;
            985: data_o = 32'h1797b7d5 /* 0x0f64 */;
            986: data_o = 32'hb7870000 /* 0x0f68 */;
            987: data_o = 32'h8e2a52a7 /* 0x0f6c */;
            988: data_o = 32'h97d38eae /* 0x0f70 */;
            989: data_o = 32'h8f32a2a7 /* 0x0f74 */;
            990: data_o = 32'h7793c78d /* 0x0f78 */;
            991: data_o = 32'hcf810048 /* 0x0f7c */;
            992: data_o = 32'h00001697 /* 0x0f80 */;
            993: data_o = 32'h27868693 /* 0x0f84 */;
            994: data_o = 32'h87ba4611 /* 0x0f88 */;
            995: data_o = 32'h873285f6 /* 0x0f8c */;
            996: data_o = 32'h867a8572 /* 0x0f90 */;
            997: data_o = 32'h1697bf55 /* 0x0f94 */;
            998: data_o = 32'h86930000 /* 0x0f98 */;
            999: data_o = 32'h460d26a6 /* 0x0f9c */;
            1000: data_o = 32'h1797b7ed /* 0x0fa0 */;
            1001: data_o = 32'hb7870000 /* 0x0fa4 */;
            1002: data_o = 32'h97d35767 /* 0x0fa8 */;
            1003: data_o = 32'heb81a2a7 /* 0x0fac */;
            1004: data_o = 32'h00001797 /* 0x0fb0 */;
            1005: data_o = 32'h5707b787 /* 0x0fb4 */;
            1006: data_o = 32'ha2f517d3 /* 0x0fb8 */;
            1007: data_o = 32'h87c2c791 /* 0x0fbc */;
            1008: data_o = 32'h85f6867a /* 0x0fc0 */;
            1009: data_o = 32'hb9558572 /* 0x0fc4 */;
            1010: data_o = 32'hf20007d3 /* 0x0fc8 */;
            1011: data_o = 32'hf4067179 /* 0x0fcc */;
            1012: data_o = 32'ha2f517d3 /* 0x0fd0 */;
            1013: data_o = 32'hc7814601 /* 0x0fd4 */;
            1014: data_o = 32'h0aa7f553 /* 0x0fd8 */;
            1015: data_o = 32'h77934605 /* 0x0fdc */;
            1016: data_o = 32'hc3c54008 /* 0x0fe0 */;
            1017: data_o = 32'h47a54881 /* 0x0fe4 */;
            1018: data_o = 32'h03000593 /* 0x0fe8 */;
            1019: data_o = 32'h02000513 /* 0x0fec */;
            1020: data_o = 32'h00d7fa63 /* 0x0ff0 */;
            1021: data_o = 32'h01110333 /* 0x0ff4 */;
            1022: data_o = 32'h00b30023 /* 0x0ff8 */;
            1023: data_o = 32'h36fd0885 /* 0x0ffc */;
            1024: data_o = 32'hfea898e3 /* 0x1000 */;
            1025: data_o = 32'hc20515d3 /* 0x1004 */;
            1026: data_o = 32'h02069f93 /* 0x1008 */;
            1027: data_o = 32'hd20587d3 /* 0x100c */;
            1028: data_o = 32'h01dfd313 /* 0x1010 */;
            1029: data_o = 32'h0a418793 /* 0x1014 */;
            1030: data_o = 32'h0af577d3 /* 0x1018 */;
            1031: data_o = 32'h2394979a /* 0x101c */;
            1032: data_o = 32'h00001797 /* 0x1020 */;
            1033: data_o = 32'h0005851b /* 0x1024 */;
            1034: data_o = 32'h12d7f7d3 /* 0x1028 */;
            1035: data_o = 32'hc2379353 /* 0x102c */;
            1036: data_o = 32'hd2337753 /* 0x1030 */;
            1037: data_o = 32'h0ae7f7d3 /* 0x1034 */;
            1038: data_o = 32'h4a87b707 /* 0x1038 */;
            1039: data_o = 32'ha2f717d3 /* 0x103c */;
            1040: data_o = 32'h0305c3b9 /* 0x1040 */;
            1041: data_o = 32'hd23377d3 /* 0x1044 */;
            1042: data_o = 32'ha2f687d3 /* 0x1048 */;
            1043: data_o = 32'h851bc781 /* 0x104c */;
            1044: data_o = 32'h43010015 /* 0x1050 */;
            1045: data_o = 32'h0f93c2b9 /* 0x1054 */;
            1046: data_o = 32'h45a90200 /* 0x1058 */;
            1047: data_o = 32'h806342a5 /* 0x105c */;
            1048: data_o = 32'h77b307f8 /* 0x1060 */;
            1049: data_o = 32'h088502b3 /* 0x1064 */;
            1050: data_o = 32'h011103b3 /* 0x1068 */;
            1051: data_o = 32'h879b36fd /* 0x106c */;
            1052: data_o = 32'h8fa30307 /* 0x1070 */;
            1053: data_o = 32'h57b3fef3 /* 0x1074 */;
            1054: data_o = 32'hfb6302b3 /* 0x1078 */;
            1055: data_o = 32'h833e0a62 /* 0x107c */;
            1056: data_o = 32'h4699bff9 /* 0x1080 */;
            1057: data_o = 32'h97d3b785 /* 0x1084 */;
            1058: data_o = 32'hf7e9a2e7 /* 0x1088 */;
            1059: data_o = 32'h00030563 /* 0x108c */;
            1060: data_o = 32'h00137793 /* 0x1090 */;
            1061: data_o = 32'h0305d3e1 /* 0x1094 */;
            1062: data_o = 32'h07d3bf75 /* 0x1098 */;
            1063: data_o = 32'h1797d205 /* 0x109c */;
            1064: data_o = 32'h75530000 /* 0x10a0 */;
            1065: data_o = 32'hb7870af5 /* 0x10a4 */;
            1066: data_o = 32'h17d342a7 /* 0x10a8 */;
            1067: data_o = 32'hc781a2f5 /* 0x10ac */;
            1068: data_o = 32'ha2a797d3 /* 0x10b0 */;
            1069: data_o = 32'h7793c789 /* 0x10b4 */;
            1070: data_o = 32'hc3910015 /* 0x10b8 */;
            1071: data_o = 32'h05932505 /* 0x10bc */;
            1072: data_o = 32'h46a90200 /* 0x10c0 */;
            1073: data_o = 32'h00b88e63 /* 0x10c4 */;
            1074: data_o = 32'h02d567bb /* 0x10c8 */;
            1075: data_o = 32'h03330885 /* 0x10cc */;
            1076: data_o = 32'h453b0111 /* 0x10d0 */;
            1077: data_o = 32'h879b02d5 /* 0x10d4 */;
            1078: data_o = 32'h0fa30307 /* 0x10d8 */;
            1079: data_o = 32'hf17dfef3 /* 0x10dc */;
            1080: data_o = 32'h00387793 /* 0x10e0 */;
            1081: data_o = 32'h94634685 /* 0x10e4 */;
            1082: data_o = 32'hc35108d7 /* 0x10e8 */;
            1083: data_o = 32'h7793e601 /* 0x10ec */;
            1084: data_o = 32'hc39100c8 /* 0x10f0 */;
            1085: data_o = 32'h1693377d /* 0x10f4 */;
            1086: data_o = 32'h92810207 /* 0x10f8 */;
            1087: data_o = 32'h02000793 /* 0x10fc */;
            1088: data_o = 32'h03000593 /* 0x1100 */;
            1089: data_o = 32'h930aa0b1 /* 0x1104 */;
            1090: data_o = 32'h01f30023 /* 0x1108 */;
            1091: data_o = 32'h09638346 /* 0x110c */;
            1092: data_o = 32'h079b02b3 /* 0x1110 */;
            1093: data_o = 32'h08930003 /* 0x1114 */;
            1094: data_o = 32'h96e30013 /* 0x1118 */;
            1095: data_o = 32'h0793fef6 /* 0x111c */;
            1096: data_o = 32'h83330203 /* 0x1120 */;
            1097: data_o = 32'h07930027 /* 0x1124 */;
            1098: data_o = 32'h002302e0 /* 0x1128 */;
            1099: data_o = 32'hbf41fef3 /* 0x112c */;
            1100: data_o = 32'h05938346 /* 0x1130 */;
            1101: data_o = 32'h86bb0200 /* 0x1134 */;
            1102: data_o = 32'h0f9300d8 /* 0x1138 */;
            1103: data_o = 32'hbfc10300 /* 0x113c */;
            1104: data_o = 32'h02000893 /* 0x1140 */;
            1105: data_o = 32'h0533bfad /* 0x1144 */;
            1106: data_o = 32'h00230111 /* 0x1148 */;
            1107: data_o = 32'h088500b5 /* 0x114c */;
            1108: data_o = 32'h00d8ff63 /* 0x1150 */;
            1109: data_o = 32'hfef899e3 /* 0x1154 */;
            1110: data_o = 32'h868a87ba /* 0x1158 */;
            1111: data_o = 32'h867a8746 /* 0x115c */;
            1112: data_o = 32'h857285f6 /* 0x1160 */;
            1113: data_o = 32'h88fff0ef /* 0x1164 */;
            1114: data_o = 32'h614570a2 /* 0x1168 */;
            1115: data_o = 32'h07938082 /* 0x116c */;
            1116: data_o = 32'h83e30200 /* 0x1170 */;
            1117: data_o = 32'hca11fef8 /* 0x1174 */;
            1118: data_o = 32'h02088793 /* 0x1178 */;
            1119: data_o = 32'h0693978a /* 0x117c */;
            1120: data_o = 32'h802302d0 /* 0x1180 */;
            1121: data_o = 32'h0885fed7 /* 0x1184 */;
            1122: data_o = 32'h7693bfc1 /* 0x1188 */;
            1123: data_o = 32'hc6990048 /* 0x118c */;
            1124: data_o = 32'h02088793 /* 0x1190 */;
            1125: data_o = 32'h0693978a /* 0x1194 */;
            1126: data_o = 32'hb7e502b0 /* 0x1198 */;
            1127: data_o = 32'h00887693 /* 0x119c */;
            1128: data_o = 32'h8693dec5 /* 0x11a0 */;
            1129: data_o = 32'h968a0208 /* 0x11a4 */;
            1130: data_o = 32'hfef68023 /* 0x11a8 */;
            1131: data_o = 32'h6783bfe9 /* 0x11ac */;
            1132: data_o = 32'h61140105 /* 0x11b0 */;
            1133: data_o = 32'h0fff0637 /* 0x11b4 */;
            1134: data_o = 32'h078a0799 /* 0x11b8 */;
            1135: data_o = 32'h439897b6 /* 0x11bc */;
            1136: data_o = 32'h93411742 /* 0x11c0 */;
            1137: data_o = 32'hc3988f51 /* 0x11c4 */;
            1138: data_o = 32'h2785491c /* 0x11c8 */;
            1139: data_o = 32'h07998b85 /* 0x11cc */;
            1140: data_o = 32'h96be078a /* 0x11d0 */;
            1141: data_o = 32'h8082c298 /* 0x11d4 */;
            1142: data_o = 32'h873e455c /* 0x11d8 */;
            1143: data_o = 32'h00f5f363 /* 0x11dc */;
            1144: data_o = 32'h451c872e /* 0x11e0 */;
            1145: data_o = 32'h0017171b /* 0x11e4 */;
            1146: data_o = 32'h17829fb9 /* 0x11e8 */;
            1147: data_o = 32'h17029381 /* 0x11ec */;
            1148: data_o = 32'h17fd9301 /* 0x11f0 */;
            1149: data_o = 32'h02e7d7b3 /* 0x11f4 */;
            1150: data_o = 32'h177d6741 /* 0x11f8 */;
            1151: data_o = 32'hf63317fd /* 0x11fc */;
            1152: data_o = 32'h836300e7 /* 0x1200 */;
            1153: data_o = 32'h863a00c7 /* 0x1204 */;
            1154: data_o = 32'h01056783 /* 0x1208 */;
            1155: data_o = 32'h75c16114 /* 0x120c */;
            1156: data_o = 32'h078a0799 /* 0x1210 */;
            1157: data_o = 32'h439897b6 /* 0x1214 */;
            1158: data_o = 32'h8f518f6d /* 0x1218 */;
            1159: data_o = 32'hc3982701 /* 0x121c */;
            1160: data_o = 32'h2785491c /* 0x1220 */;
            1161: data_o = 32'h07998b85 /* 0x1224 */;
            1162: data_o = 32'h96be078a /* 0x1228 */;
            1163: data_o = 32'h8082c298 /* 0x122c */;
            1164: data_o = 32'h0737611c /* 0x1230 */;
            1165: data_o = 32'h46374000 /* 0x1234 */;
            1166: data_o = 32'ha223000f /* 0x1238 */;
            1167: data_o = 32'haa230007 /* 0x123c */;
            1168: data_o = 32'hcb980207 /* 0x1240 */;
            1169: data_o = 32'h24060613 /* 0x1244 */;
            1170: data_o = 32'h400005b7 /* 0x1248 */;
            1171: data_o = 32'h367d4bd8 /* 0x124c */;
            1172: data_o = 32'he6012701 /* 0x1250 */;
            1173: data_o = 32'h0007a823 /* 0x1254 */;
            1174: data_o = 32'h76b38082 /* 0x1258 */;
            1175: data_o = 32'h171b00b7 /* 0x125c */;
            1176: data_o = 32'h8f550107 /* 0x1260 */;
            1177: data_o = 32'hf37d2701 /* 0x1264 */;
            1178: data_o = 32'h80000737 /* 0x1268 */;
            1179: data_o = 32'h4918cb98 /* 0x126c */;
            1180: data_o = 32'h8b052705 /* 0x1270 */;
            1181: data_o = 32'h4bdcd398 /* 0x1274 */;
            1182: data_o = 32'h0167d79b /* 0x1278 */;
            1183: data_o = 32'h0c238b85 /* 0x127c */;
            1184: data_o = 32'h808200f5 /* 0x1280 */;
            1185: data_o = 32'h02069713 /* 0x1284 */;
            1186: data_o = 32'h19c18793 /* 0x1288 */;
            1187: data_o = 32'h71599301 /* 0x128c */;
            1188: data_o = 32'hf0a297ba /* 0x1290 */;
            1189: data_o = 32'h0007c403 /* 0x1294 */;
            1190: data_o = 32'hf486e4ce /* 0x1298 */;
            1191: data_o = 32'h0034099b /* 0x129c */;
            1192: data_o = 32'he8caeca6 /* 0x12a0 */;
            1193: data_o = 32'hfc56e0d2 /* 0x12a4 */;
            1194: data_o = 32'hf45ef85a /* 0x12a8 */;
            1195: data_o = 32'hec66f062 /* 0x12ac */;
            1196: data_o = 32'hf993e86a /* 0x12b0 */;
            1197: data_o = 32'h47a11fc9 /* 0x12b4 */;
            1198: data_o = 32'h1337e063 /* 0x12b8 */;
            1199: data_o = 32'h0285d793 /* 0x12bc */;
            1200: data_o = 32'h00f10023 /* 0x12c0 */;
            1201: data_o = 32'h0205d793 /* 0x12c4 */;
            1202: data_o = 32'h00f100a3 /* 0x12c8 */;
            1203: data_o = 32'h0105d793 /* 0x12cc */;
            1204: data_o = 32'h00f101a3 /* 0x12d0 */;
            1205: data_o = 32'h0085979b /* 0x12d4 */;
            1206: data_o = 32'h0105959b /* 0x12d8 */;
            1207: data_o = 32'h0105d59b /* 0x12dc */;
            1208: data_o = 32'h0085d59b /* 0x12e0 */;
            1209: data_o = 32'h8a328fcd /* 0x12e4 */;
            1210: data_o = 32'h47058936 /* 0x12e8 */;
            1211: data_o = 32'h860a4681 /* 0x12ec */;
            1212: data_o = 32'h03000593 /* 0x12f0 */;
            1213: data_o = 32'h012384aa /* 0x12f4 */;
            1214: data_o = 32'h12230001 /* 0x12f8 */;
            1215: data_o = 32'he0ef00f1 /* 0x12fc */;
            1216: data_o = 32'hed21f93f /* 0x1300 */;
            1217: data_o = 32'h9c132401 /* 0x1304 */;
            1218: data_o = 32'h4b810039 /* 0x1308 */;
            1219: data_o = 32'h4b014a85 /* 0x130c */;
            1220: data_o = 32'h0d134c85 /* 0x1310 */;
            1221: data_o = 32'he02504c0 /* 0x1314 */;
            1222: data_o = 32'h1b634785 /* 0x1318 */;
            1223: data_o = 32'h896302f9 /* 0x131c */;
            1224: data_o = 32'h6409020a /* 0x1320 */;
            1225: data_o = 32'h71040413 /* 0x1324 */;
            1226: data_o = 32'h47014911 /* 0x1328 */;
            1227: data_o = 32'h46010034 /* 0x132c */;
            1228: data_o = 32'h02000593 /* 0x1330 */;
            1229: data_o = 32'hf0ef8526 /* 0x1334 */;
            1230: data_o = 32'h4781af0f /* 0x1338 */;
            1231: data_o = 32'h973e0038 /* 0x133c */;
            1232: data_o = 32'h00074703 /* 0x1340 */;
            1233: data_o = 32'h0785e711 /* 0x1344 */;
            1234: data_o = 32'hff279ae3 /* 0x1348 */;
            1235: data_o = 32'hfc71347d /* 0x134c */;
            1236: data_o = 32'h45814609 /* 0x1350 */;
            1237: data_o = 32'he0ef8526 /* 0x1354 */;
            1238: data_o = 32'h70a6ea9f /* 0x1358 */;
            1239: data_o = 32'h64e67406 /* 0x135c */;
            1240: data_o = 32'h69a66946 /* 0x1360 */;
            1241: data_o = 32'h7ae26a06 /* 0x1364 */;
            1242: data_o = 32'h7ba27b42 /* 0x1368 */;
            1243: data_o = 32'h6ce27c02 /* 0x136c */;
            1244: data_o = 32'h61656d42 /* 0x1370 */;
            1245: data_o = 32'h47018082 /* 0x1374 */;
            1246: data_o = 32'h46010034 /* 0x1378 */;
            1247: data_o = 32'h852685e2 /* 0x137c */;
            1248: data_o = 32'haa6ff0ef /* 0x1380 */;
            1249: data_o = 32'h4683f979 /* 0x1384 */;
            1250: data_o = 32'h003c0001 /* 0x1388 */;
            1251: data_o = 32'h84e34701 /* 0x138c */;
            1252: data_o = 32'h9463f8e9 /* 0x1390 */;
            1253: data_o = 32'h8f63000b /* 0x1394 */;
            1254: data_o = 32'h166303a6 /* 0x1398 */;
            1255: data_o = 32'h8603000b /* 0x139c */;
            1256: data_o = 32'h4b630007 /* 0x13a0 */;
            1257: data_o = 32'hcc010006 /* 0x13a4 */;
            1258: data_o = 32'h0007c583 /* 0x13a8 */;
            1259: data_o = 32'h008a0633 /* 0x13ac */;
            1260: data_o = 32'h0fa34b05 /* 0x13b0 */;
            1261: data_o = 32'h347dfeb6 /* 0x13b4 */;
            1262: data_o = 32'h07852705 /* 0x13b8 */;
            1263: data_o = 32'h4b05bfc9 /* 0x13bc */;
            1264: data_o = 32'hff991ce3 /* 0x13c0 */;
            1265: data_o = 32'hfe0a8ae3 /* 0x13c4 */;
            1266: data_o = 32'h0007c603 /* 0x13c8 */;
            1267: data_o = 32'h3a938b56 /* 0x13cc */;
            1268: data_o = 32'hb7dd0016 /* 0x13d0 */;
            1269: data_o = 32'hb7cd4b85 /* 0x13d4 */;
            1270: data_o = 32'hb741557d /* 0x13d8 */;
            1271: data_o = 32'h971b7175 /* 0x13dc */;
            1272: data_o = 32'he1220085 /* 0x13e0 */;
            1273: data_o = 32'hf8cafca6 /* 0x13e4 */;
            1274: data_o = 32'he5061702 /* 0x13e8 */;
            1275: data_o = 32'hf0d2f4ce /* 0x13ec */;
            1276: data_o = 32'he8daecd6 /* 0x13f0 */;
            1277: data_o = 32'he0e2e4de /* 0x13f4 */;
            1278: data_o = 32'hf86afc66 /* 0x13f8 */;
            1279: data_o = 32'h4785f46e /* 0x13fc */;
            1280: data_o = 32'h84b2892a /* 0x1400 */;
            1281: data_o = 32'h93018436 /* 0x1404 */;
            1282: data_o = 32'h0cf69963 /* 0x1408 */;
            1283: data_o = 32'h05100793 /* 0x140c */;
            1284: data_o = 32'h8f5d17a2 /* 0x1410 */;
            1285: data_o = 32'h579be83a /* 0x1414 */;
            1286: data_o = 32'h46810187 /* 0x1418 */;
            1287: data_o = 32'h45894601 /* 0x141c */;
            1288: data_o = 32'h02800813 /* 0x1420 */;
            1289: data_o = 32'hd51348a1 /* 0x1424 */;
            1290: data_o = 32'hcd4500f7 /* 0x1428 */;
            1291: data_o = 32'h05137565 /* 0x142c */;
            1292: data_o = 32'h08139005 /* 0x1430 */;
            1293: data_o = 32'h08930270 /* 0x1434 */;
            1294: data_o = 32'h43210280 /* 0x1438 */;
            1295: data_o = 32'h17c28fa9 /* 0x143c */;
            1296: data_o = 32'hde1393c1 /* 0x1440 */;
            1297: data_o = 32'h186300f7 /* 0x1444 */;
            1298: data_o = 32'h71630e0e /* 0x1448 */;
            1299: data_o = 32'hd79b0cd8 /* 0x144c */;
            1300: data_o = 32'h979b0097 /* 0x1450 */;
            1301: data_o = 32'hd79b0107 /* 0x1454 */;
            1302: data_o = 32'h979b0107 /* 0x1458 */;
            1303: data_o = 32'he7930017 /* 0x145c */;
            1304: data_o = 32'h27810017 /* 0x1460 */;
            1305: data_o = 32'hd7138fd9 /* 0x1464 */;
            1306: data_o = 32'h04230287 /* 0x1468 */;
            1307: data_o = 32'hd71300e1 /* 0x146c */;
            1308: data_o = 32'h05230187 /* 0x1470 */;
            1309: data_o = 32'hd71300e1 /* 0x1474 */;
            1310: data_o = 32'he83e0107 /* 0x1478 */;
            1311: data_o = 32'h00e105a3 /* 0x147c */;
            1312: data_o = 32'h0087971b /* 0x1480 */;
            1313: data_o = 32'h0107979b /* 0x1484 */;
            1314: data_o = 32'h0107d79b /* 0x1488 */;
            1315: data_o = 32'h0087d79b /* 0x148c */;
            1316: data_o = 32'h46818fd9 /* 0x1490 */;
            1317: data_o = 32'h00304705 /* 0x1494 */;
            1318: data_o = 32'h03000593 /* 0x1498 */;
            1319: data_o = 32'h04a3854a /* 0x149c */;
            1320: data_o = 32'h16230001 /* 0x14a0 */;
            1321: data_o = 32'he0ef00f1 /* 0x14a4 */;
            1322: data_o = 32'h89aadebf /* 0x14a8 */;
            1323: data_o = 32'h1a051663 /* 0x14ac */;
            1324: data_o = 32'h4a814a01 /* 0x14b0 */;
            1325: data_o = 32'h0fe00b13 /* 0x14b4 */;
            1326: data_o = 32'h11634b91 /* 0x14b8 */;
            1327: data_o = 32'h47850944 /* 0x14bc */;
            1328: data_o = 32'h22f40463 /* 0x14c0 */;
            1329: data_o = 32'h15aa45cd /* 0x14c4 */;
            1330: data_o = 32'h08304685 /* 0x14c8 */;
            1331: data_o = 32'h06158593 /* 0x14cc */;
            1332: data_o = 32'hec02854a /* 0x14d0 */;
            1333: data_o = 32'hdb1ff0ef /* 0x14d4 */;
            1334: data_o = 32'h0793aabd /* 0x14d8 */;
            1335: data_o = 32'h17a60290 /* 0x14dc */;
            1336: data_o = 32'h979bbf0d /* 0x14e0 */;
            1337: data_o = 32'h17c20017 /* 0x14e4 */;
            1338: data_o = 32'h93c12685 /* 0x14e8 */;
            1339: data_o = 32'h80e32605 /* 0x14ec */;
            1340: data_o = 32'h1ae3f706 /* 0x14f0 */;
            1341: data_o = 32'h58e3f316 /* 0x14f4 */;
            1342: data_o = 32'h8613f2b0 /* 0x14f8 */;
            1343: data_o = 32'h960a0205 /* 0x14fc */;
            1344: data_o = 32'hff064603 /* 0x1500 */;
            1345: data_o = 32'h8fd135fd /* 0x1504 */;
            1346: data_o = 32'hbf314601 /* 0x1508 */;
            1347: data_o = 32'h0017979b /* 0x150c */;
            1348: data_o = 32'h268517c2 /* 0x1510 */;
            1349: data_o = 32'h260593c1 /* 0x1514 */;
            1350: data_o = 32'hf3168be3 /* 0x1518 */;
            1351: data_o = 32'hf26613e3 /* 0x151c */;
            1352: data_o = 32'hf2b051e3 /* 0x1520 */;
            1353: data_o = 32'h02058613 /* 0x1524 */;
            1354: data_o = 32'h4603960a /* 0x1528 */;
            1355: data_o = 32'h35fdff06 /* 0x152c */;
            1356: data_o = 32'h46018fd1 /* 0x1530 */;
            1357: data_o = 32'h73e3b739 /* 0x1534 */;
            1358: data_o = 32'hbf11f0d8 /* 0x1538 */;
            1359: data_o = 32'h1c1b2a05 /* 0x153c */;
            1360: data_o = 32'h0d9b009a /* 0x1540 */;
            1361: data_o = 32'h0d13000c /* 0x1544 */;
            1362: data_o = 32'h47012000 /* 0x1548 */;
            1363: data_o = 32'h46010834 /* 0x154c */;
            1364: data_o = 32'h02000593 /* 0x1550 */;
            1365: data_o = 32'he0ef854a /* 0x1554 */;
            1366: data_o = 32'h1e63d3bf /* 0x1558 */;
            1367: data_o = 32'h08300e05 /* 0x155c */;
            1368: data_o = 32'h46814c81 /* 0x1560 */;
            1369: data_o = 32'h00064783 /* 0x1564 */;
            1370: data_o = 32'h10069863 /* 0x1568 */;
            1371: data_o = 32'h0c0a9363 /* 0x156c */;
            1372: data_o = 32'hca93839d /* 0x1570 */;
            1373: data_o = 32'h2c850017 /* 0x1574 */;
            1374: data_o = 32'h95e30605 /* 0x1578 */;
            1375: data_o = 32'hd6f1ff7c /* 0x157c */;
            1376: data_o = 32'h020c1693 /* 0x1580 */;
            1377: data_o = 32'h020d1793 /* 0x1584 */;
            1378: data_o = 32'h93819281 /* 0x1588 */;
            1379: data_o = 32'h159b8e9d /* 0x158c */;
            1380: data_o = 32'h4701003d /* 0x1590 */;
            1381: data_o = 32'h460196a6 /* 0x1594 */;
            1382: data_o = 32'hf0ef854a /* 0x1598 */;
            1383: data_o = 32'hed4588cf /* 0x159c */;
            1384: data_o = 32'h08344701 /* 0x15a0 */;
            1385: data_o = 32'h45c14601 /* 0x15a4 */;
            1386: data_o = 32'he0ef854a /* 0x15a8 */;
            1387: data_o = 32'he545ce7f /* 0x15ac */;
            1388: data_o = 32'h01815683 /* 0x15b0 */;
            1389: data_o = 32'he00c0c1b /* 0x15b4 */;
            1390: data_o = 32'h5c131c02 /* 0x15b8 */;
            1391: data_o = 32'h9c26020c /* 0x15bc */;
            1392: data_o = 32'h0086979b /* 0x15c0 */;
            1393: data_o = 32'h8edd82a1 /* 0x15c4 */;
            1394: data_o = 32'h000c4703 /* 0x15c8 */;
            1395: data_o = 32'h001c4783 /* 0x15cc */;
            1396: data_o = 32'h0106969b /* 0x15d0 */;
            1397: data_o = 32'h0187171b /* 0x15d4 */;
            1398: data_o = 32'h0107979b /* 0x15d8 */;
            1399: data_o = 32'h47038fd9 /* 0x15dc */;
            1400: data_o = 32'hd69b003c /* 0x15e0 */;
            1401: data_o = 32'h46014106 /* 0x15e4 */;
            1402: data_o = 32'h47038fd9 /* 0x15e8 */;
            1403: data_o = 32'h6505002c /* 0x15ec */;
            1404: data_o = 32'h171b4821 /* 0x15f0 */;
            1405: data_o = 32'h8fd90087 /* 0x15f4 */;
            1406: data_o = 32'h47012781 /* 0x15f8 */;
            1407: data_o = 32'h1ff00893 /* 0x15fc */;
            1408: data_o = 32'h0807d763 /* 0x1600 */;
            1409: data_o = 32'h88108837 /* 0x1604 */;
            1410: data_o = 32'h48a16585 /* 0x1608 */;
            1411: data_o = 32'h1ff00313 /* 0x160c */;
            1412: data_o = 32'h0107c7b3 /* 0x1610 */;
            1413: data_o = 32'hc6632781 /* 0x1614 */;
            1414: data_o = 32'h6f630c07 /* 0x1618 */;
            1415: data_o = 32'hd79b08b6 /* 0x161c */;
            1416: data_o = 32'h979b0107 /* 0x1620 */;
            1417: data_o = 32'hd79b0107 /* 0x1624 */;
            1418: data_o = 32'h88e34107 /* 0x1628 */;
            1419: data_o = 32'h557de8d7 /* 0x162c */;
            1420: data_o = 32'h8c63a01d /* 0x1630 */;
            1421: data_o = 32'hf7930567 /* 0x1634 */;
            1422: data_o = 32'hff950f07 /* 0x1638 */;
            1423: data_o = 32'h46814709 /* 0x163c */;
            1424: data_o = 32'h45814601 /* 0x1640 */;
            1425: data_o = 32'he0ef854a /* 0x1644 */;
            1426: data_o = 32'h8793fe1f /* 0x1648 */;
            1427: data_o = 32'h8cb3020c /* 0x164c */;
            1428: data_o = 32'hc5030027 /* 0x1650 */;
            1429: data_o = 32'h89aaff8c /* 0x1654 */;
            1430: data_o = 32'h640a60aa /* 0x1658 */;
            1431: data_o = 32'h794674e6 /* 0x165c */;
            1432: data_o = 32'h6ae67a06 /* 0x1660 */;
            1433: data_o = 32'h6ba66b46 /* 0x1664 */;
            1434: data_o = 32'h7ce26c06 /* 0x1668 */;
            1435: data_o = 32'h7da27d42 /* 0x166c */;
            1436: data_o = 32'h79a6854e /* 0x1670 */;
            1437: data_o = 32'h80826149 /* 0x1674 */;
            1438: data_o = 32'h41ad873b /* 0x1678 */;
            1439: data_o = 32'h93011702 /* 0x167c */;
            1440: data_o = 32'h00239726 /* 0x1680 */;
            1441: data_o = 32'h3d7d00f7 /* 0x1684 */;
            1442: data_o = 32'h86d6b5fd /* 0x1688 */;
            1443: data_o = 32'h959bb5ed /* 0x168c */;
            1444: data_o = 32'h26050017 /* 0x1690 */;
            1445: data_o = 32'h0005879b /* 0x1694 */;
            1446: data_o = 32'h02e32705 /* 0x1698 */;
            1447: data_o = 32'h11e3f8a6 /* 0x169c */;
            1448: data_o = 32'hcfe3f707 /* 0x16a0 */;
            1449: data_o = 32'h07b3f598 /* 0x16a4 */;
            1450: data_o = 32'hc783019c /* 0x16a8 */;
            1451: data_o = 32'h2c850007 /* 0x16ac */;
            1452: data_o = 32'h8fcd4701 /* 0x16b0 */;
            1453: data_o = 32'hb7a92781 /* 0x16b4 */;
            1454: data_o = 32'h0017951b /* 0x16b8 */;
            1455: data_o = 32'h079b2605 /* 0x16bc */;
            1456: data_o = 32'h27050005 /* 0x16c0 */;
            1457: data_o = 32'hf4b60de3 /* 0x16c4 */;
            1458: data_o = 32'hf51717e3 /* 0x16c8 */;
            1459: data_o = 32'hf59345e3 /* 0x16cc */;
            1460: data_o = 32'h019c07b3 /* 0x16d0 */;
            1461: data_o = 32'h0007c783 /* 0x16d4 */;
            1462: data_o = 32'h47012c85 /* 0x16d8 */;
            1463: data_o = 32'h27818fc9 /* 0x16dc */;
            1464: data_o = 32'h67e3bf1d /* 0x16e0 */;
            1465: data_o = 32'hbf25f2b6 /* 0x16e4 */;
            1466: data_o = 32'h46814709 /* 0x16e8 */;
            1467: data_o = 32'h45814601 /* 0x16ec */;
            1468: data_o = 32'he0ef854a /* 0x16f0 */;
            1469: data_o = 32'hb78df35f /* 0x16f4 */;
            1470: data_o = 32'hb1cdc291 /* 0x16f8 */;
            1471: data_o = 32'h80824501 /* 0x16fc */;
            1472: data_o = 32'hf1227151 /* 0x1700 */;
            1473: data_o = 32'he152e54e /* 0x1704 */;
            1474: data_o = 32'h1920fcd6 /* 0x1708 */;
            1475: data_o = 32'h6a2569c1 /* 0x170c */;
            1476: data_o = 32'hed266a85 /* 0x1710 */;
            1477: data_o = 32'hf8dae94a /* 0x1714 */;
            1478: data_o = 32'hf4def506 /* 0x1718 */;
            1479: data_o = 32'hece6f0e2 /* 0x171c */;
            1480: data_o = 32'he4eee8ea /* 0x1720 */;
            1481: data_o = 32'hfd2e892a /* 0x1724 */;
            1482: data_o = 32'he5b6e1b2 /* 0x1728 */;
            1483: data_o = 32'hedbee9ba /* 0x172c */;
            1484: data_o = 32'hf5c6f1c2 /* 0x1730 */;
            1485: data_o = 32'h4481fc22 /* 0x1734 */;
            1486: data_o = 32'h02500b13 /* 0x1738 */;
            1487: data_o = 32'h0a1319fd /* 0x173c */;
            1488: data_o = 32'h8a93041a /* 0x1740 */;
            1489: data_o = 32'h4503800a /* 0x1744 */;
            1490: data_o = 32'hed050009 /* 0x1748 */;
            1491: data_o = 32'h862657f9 /* 0x174c */;
            1492: data_o = 32'h0097f363 /* 0x1750 */;
            1493: data_o = 32'h180c5679 /* 0x1754 */;
            1494: data_o = 32'h56fd4501 /* 0x1758 */;
            1495: data_o = 32'ha85fe0ef /* 0x175c */;
            1496: data_o = 32'h740a70aa /* 0x1760 */;
            1497: data_o = 32'h69aa694a /* 0x1764 */;
            1498: data_o = 32'h7ae66a0a /* 0x1768 */;
            1499: data_o = 32'h7ba67b46 /* 0x176c */;
            1500: data_o = 32'h6ce67c06 /* 0x1770 */;
            1501: data_o = 32'h6da66d46 /* 0x1774 */;
            1502: data_o = 32'h0004851b /* 0x1778 */;
            1503: data_o = 32'h616d64ea /* 0x177c */;
            1504: data_o = 32'h09058082 /* 0x1780 */;
            1505: data_o = 32'h01650863 /* 0x1784 */;
            1506: data_o = 32'h00148b93 /* 0x1788 */;
            1507: data_o = 32'h862656fd /* 0x178c */;
            1508: data_o = 32'haabd180c /* 0x1790 */;
            1509: data_o = 32'h07134581 /* 0x1794 */;
            1510: data_o = 32'h061302b0 /* 0x1798 */;
            1511: data_o = 32'h051302d0 /* 0x179c */;
            1512: data_o = 32'h08130300 /* 0x17a0 */;
            1513: data_o = 32'h08930200 /* 0x17a4 */;
            1514: data_o = 32'ha8010230 /* 0x17a8 */;
            1515: data_o = 32'h02c78e63 /* 0x17ac */;
            1516: data_o = 32'h02a79163 /* 0x17b0 */;
            1517: data_o = 32'h0015e593 /* 0x17b4 */;
            1518: data_o = 32'h47838936 /* 0x17b8 */;
            1519: data_o = 32'h06930009 /* 0x17bc */;
            1520: data_o = 32'h86630019 /* 0x17c0 */;
            1521: data_o = 32'h63e302e7 /* 0x17c4 */;
            1522: data_o = 32'h8563fef7 /* 0x17c8 */;
            1523: data_o = 32'h86630307 /* 0x17cc */;
            1524: data_o = 32'h871b0317 /* 0x17d0 */;
            1525: data_o = 32'h7713fd07 /* 0x17d4 */;
            1526: data_o = 32'h46250ff7 /* 0x17d8 */;
            1527: data_o = 32'h06e66a63 /* 0x17dc */;
            1528: data_o = 32'h46a54881 /* 0x17e0 */;
            1529: data_o = 32'ha0254529 /* 0x17e4 */;
            1530: data_o = 32'h0025e593 /* 0x17e8 */;
            1531: data_o = 32'he593b7f1 /* 0x17ec */;
            1532: data_o = 32'hb7d90045 /* 0x17f0 */;
            1533: data_o = 32'h0085e593 /* 0x17f4 */;
            1534: data_o = 32'he593b7c1 /* 0x17f8 */;
            1535: data_o = 32'hbf6d0105 /* 0x17fc */;
            1536: data_o = 32'h031508bb /* 0x1800 */;
            1537: data_o = 32'h889b8932 /* 0x1804 */;
            1538: data_o = 32'h88bbfd08 /* 0x1808 */;
            1539: data_o = 32'h470300e8 /* 0x180c */;
            1540: data_o = 32'h06130009 /* 0x1810 */;
            1541: data_o = 32'h079b0019 /* 0x1814 */;
            1542: data_o = 32'hf793fd07 /* 0x1818 */;
            1543: data_o = 32'hf1e30ff7 /* 0x181c */;
            1544: data_o = 32'h4703fef6 /* 0x1820 */;
            1545: data_o = 32'h07930009 /* 0x1824 */;
            1546: data_o = 32'h480102e0 /* 0x1828 */;
            1547: data_o = 32'h08f71663 /* 0x182c */;
            1548: data_o = 32'h00194683 /* 0x1830 */;
            1549: data_o = 32'h07934625 /* 0x1834 */;
            1550: data_o = 32'h871b0019 /* 0x1838 */;
            1551: data_o = 32'h7713fd06 /* 0x183c */;
            1552: data_o = 32'he5930ff7 /* 0x1840 */;
            1553: data_o = 32'h6b634005 /* 0x1844 */;
            1554: data_o = 32'h462504e6 /* 0x1848 */;
            1555: data_o = 32'ha81d4329 /* 0x184c */;
            1556: data_o = 32'h02a00713 /* 0x1850 */;
            1557: data_o = 32'h96e34881 /* 0x1854 */;
            1558: data_o = 32'h401cfce7 /* 0x1858 */;
            1559: data_o = 32'h00840713 /* 0x185c */;
            1560: data_o = 32'h0007889b /* 0x1860 */;
            1561: data_o = 32'h0007d663 /* 0x1864 */;
            1562: data_o = 32'h0025e593 /* 0x1868 */;
            1563: data_o = 32'h40f008bb /* 0x186c */;
            1564: data_o = 32'h8936843a /* 0x1870 */;
            1565: data_o = 32'h083bb77d /* 0x1874 */;
            1566: data_o = 32'h87aa0303 /* 0x1878 */;
            1567: data_o = 32'hfd08081b /* 0x187c */;
            1568: data_o = 32'h00d8083b /* 0x1880 */;
            1569: data_o = 32'h0007c683 /* 0x1884 */;
            1570: data_o = 32'h00178513 /* 0x1888 */;
            1571: data_o = 32'hfd06871b /* 0x188c */;
            1572: data_o = 32'h0ff77713 /* 0x1890 */;
            1573: data_o = 32'hfee671e3 /* 0x1894 */;
            1574: data_o = 32'ha839893e /* 0x1898 */;
            1575: data_o = 32'h02a00713 /* 0x189c */;
            1576: data_o = 32'hfee69ce3 /* 0x18a0 */;
            1577: data_o = 32'h0713401c /* 0x18a4 */;
            1578: data_o = 32'h881b0084 /* 0x18a8 */;
            1579: data_o = 32'hd3630007 /* 0x18ac */;
            1580: data_o = 32'h48010007 /* 0x18b0 */;
            1581: data_o = 32'h843a0909 /* 0x18b4 */;
            1582: data_o = 32'h00094783 /* 0x18b8 */;
            1583: data_o = 32'h06c00693 /* 0x18bc */;
            1584: data_o = 32'h00190713 /* 0x18c0 */;
            1585: data_o = 32'h06d78163 /* 0x18c4 */;
            1586: data_o = 32'h04f6e863 /* 0x18c8 */;
            1587: data_o = 32'h06800693 /* 0x18cc */;
            1588: data_o = 32'h06d78663 /* 0x18d0 */;
            1589: data_o = 32'h06a00693 /* 0x18d4 */;
            1590: data_o = 32'h04d78b63 /* 0x18d8 */;
            1591: data_o = 32'h00094503 /* 0x18dc */;
            1592: data_o = 32'h06700793 /* 0x18e0 */;
            1593: data_o = 32'heb630905 /* 0x18e4 */;
            1594: data_o = 32'h07930ca7 /* 0x18e8 */;
            1595: data_o = 32'he2630570 /* 0x18ec */;
            1596: data_o = 32'h079306a7 /* 0x18f0 */;
            1597: data_o = 32'h04630450 /* 0x18f4 */;
            1598: data_o = 32'hea6308f5 /* 0x18f8 */;
            1599: data_o = 32'h15e306a7 /* 0x18fc */;
            1600: data_o = 32'h8b93e965 /* 0x1900 */;
            1601: data_o = 32'h56fd0014 /* 0x1904 */;
            1602: data_o = 32'h180c8626 /* 0x1908 */;
            1603: data_o = 32'h02500513 /* 0x190c */;
            1604: data_o = 32'h8d1fe0ef /* 0x1910 */;
            1605: data_o = 32'hbd0584de /* 0x1914 */;
            1606: data_o = 32'h07400693 /* 0x1918 */;
            1607: data_o = 32'h00d78963 /* 0x191c */;
            1608: data_o = 32'h07a00693 /* 0x1920 */;
            1609: data_o = 32'h4683bf55 /* 0x1924 */;
            1610: data_o = 32'h85630019 /* 0x1928 */;
            1611: data_o = 32'he59300f6 /* 0x192c */;
            1612: data_o = 32'ha8191005 /* 0x1930 */;
            1613: data_o = 32'h3005e593 /* 0x1934 */;
            1614: data_o = 32'hb74d0909 /* 0x1938 */;
            1615: data_o = 32'h00194683 /* 0x193c */;
            1616: data_o = 32'h00f68663 /* 0x1940 */;
            1617: data_o = 32'h0805e593 /* 0x1944 */;
            1618: data_o = 32'hbf49893a /* 0x1948 */;
            1619: data_o = 32'h0c05e593 /* 0x194c */;
            1620: data_o = 32'h079bb7e5 /* 0x1950 */;
            1621: data_o = 32'hf793fa85 /* 0x1954 */;
            1622: data_o = 32'h473d0ff7 /* 0x1958 */;
            1623: data_o = 32'he2f766e3 /* 0x195c */;
            1624: data_o = 32'he7c18713 /* 0x1960 */;
            1625: data_o = 32'h97ba078a /* 0x1964 */;
            1626: data_o = 32'h97ba439c /* 0x1968 */;
            1627: data_o = 32'h07938782 /* 0x196c */;
            1628: data_o = 32'h03630460 /* 0x1970 */;
            1629: data_o = 32'h07931ef5 /* 0x1974 */;
            1630: data_o = 32'h17e30470 /* 0x1978 */;
            1631: data_o = 32'h7793e0f5 /* 0x197c */;
            1632: data_o = 32'h07130df5 /* 0x1980 */;
            1633: data_o = 32'h96630470 /* 0x1984 */;
            1634: data_o = 32'he5b300e7 /* 0x1988 */;
            1635: data_o = 32'h75130155 /* 0x198c */;
            1636: data_o = 32'h07930fd5 /* 0x1990 */;
            1637: data_o = 32'h14630450 /* 0x1994 */;
            1638: data_o = 32'he59300f5 /* 0x1998 */;
            1639: data_o = 32'h20080205 /* 0x199c */;
            1640: data_o = 32'hfffff517 /* 0x19a0 */;
            1641: data_o = 32'h874687ae /* 0x19a4 */;
            1642: data_o = 32'h862686c2 /* 0x19a8 */;
            1643: data_o = 32'h0513180c /* 0x19ac */;
            1644: data_o = 32'h0b938405 /* 0x19b0 */;
            1645: data_o = 32'hf0ef0084 /* 0x19b4 */;
            1646: data_o = 32'ha8d9ac4f /* 0x19b8 */;
            1647: data_o = 32'hf975079b /* 0x19bc */;
            1648: data_o = 32'h0ff7f793 /* 0x19c0 */;
            1649: data_o = 32'h61e3473d /* 0x19c4 */;
            1650: data_o = 32'h4705dcf7 /* 0x19c8 */;
            1651: data_o = 32'h00f71733 /* 0x19cc */;
            1652: data_o = 32'h01477733 /* 0x19d0 */;
            1653: data_o = 32'h4729e71d /* 0x19d4 */;
            1654: data_o = 32'h24e78063 /* 0x19d8 */;
            1655: data_o = 32'h95e3471d /* 0x19dc */;
            1656: data_o = 32'he593dae7 /* 0x19e0 */;
            1657: data_o = 32'he5170215 /* 0x19e4 */;
            1658: data_o = 32'h6014ffff /* 0x19e8 */;
            1659: data_o = 32'h00840b93 /* 0x19ec */;
            1660: data_o = 32'h48c1e02e /* 0x19f0 */;
            1661: data_o = 32'h470147c1 /* 0x19f4 */;
            1662: data_o = 32'h180c8626 /* 0x19f8 */;
            1663: data_o = 32'h7fa50513 /* 0x19fc */;
            1664: data_o = 32'h0713a071 /* 0x1a00 */;
            1665: data_o = 32'h47c10780 /* 0x1a04 */;
            1666: data_o = 32'h02e50863 /* 0x1a08 */;
            1667: data_o = 32'h06200793 /* 0x1a0c */;
            1668: data_o = 32'h02f50663 /* 0x1a10 */;
            1669: data_o = 32'h06f00793 /* 0x1a14 */;
            1670: data_o = 32'h30f50563 /* 0x1a18 */;
            1671: data_o = 32'h05800793 /* 0x1a1c */;
            1672: data_o = 32'h00f50963 /* 0x1a20 */;
            1673: data_o = 32'h47a999bd /* 0x1a24 */;
            1674: data_o = 32'h06900713 /* 0x1a28 */;
            1675: data_o = 32'h00e50d63 /* 0x1a2c */;
            1676: data_o = 32'he593a039 /* 0x1a30 */;
            1677: data_o = 32'h47c10205 /* 0x1a34 */;
            1678: data_o = 32'ha03199cd /* 0x1a38 */;
            1679: data_o = 32'h07134789 /* 0x1a3c */;
            1680: data_o = 32'h1be30640 /* 0x1a40 */;
            1681: data_o = 32'hf713fee5 /* 0x1a44 */;
            1682: data_o = 32'hc3114005 /* 0x1a48 */;
            1683: data_o = 32'h178299f9 /* 0x1a4c */;
            1684: data_o = 32'h06900613 /* 0x1a50 */;
            1685: data_o = 32'hf693872e /* 0x1a54 */;
            1686: data_o = 32'h93812005 /* 0x1a58 */;
            1687: data_o = 32'h00840b93 /* 0x1a5c */;
            1688: data_o = 32'h00c50663 /* 0x1a60 */;
            1689: data_o = 32'h06400613 /* 0x1a64 */;
            1690: data_o = 32'h08c51963 /* 0x1a68 */;
            1691: data_o = 32'h6018c68d /* 0x1a6c */;
            1692: data_o = 32'hffffe517 /* 0x1a70 */;
            1693: data_o = 32'h5693e02e /* 0x1a74 */;
            1694: data_o = 32'hc63343f7 /* 0x1a78 */;
            1695: data_o = 32'h06b300e6 /* 0x1a7c */;
            1696: data_o = 32'h937d40d6 /* 0x1a80 */;
            1697: data_o = 32'h180c8626 /* 0x1a84 */;
            1698: data_o = 32'h77050513 /* 0x1a88 */;
            1699: data_o = 32'h826ff0ef /* 0x1a8c */;
            1700: data_o = 32'h845e84aa /* 0x1a90 */;
            1701: data_o = 32'hf713b94d /* 0x1a94 */;
            1702: data_o = 32'h86ae1005 /* 0x1a98 */;
            1703: data_o = 32'h6018c30d /* 0x1a9c */;
            1704: data_o = 32'hffffe517 /* 0x1aa0 */;
            1705: data_o = 32'h5693e02e /* 0x1aa4 */;
            1706: data_o = 32'hc63343f7 /* 0x1aa8 */;
            1707: data_o = 32'h06b300e6 /* 0x1aac */;
            1708: data_o = 32'h937d40d6 /* 0x1ab0 */;
            1709: data_o = 32'h180c8626 /* 0x1ab4 */;
            1710: data_o = 32'h74050513 /* 0x1ab8 */;
            1711: data_o = 32'hf613bfc1 /* 0x1abc */;
            1712: data_o = 32'h40180405 /* 0x1ac0 */;
            1713: data_o = 32'h7713c21d /* 0x1ac4 */;
            1714: data_o = 32'h569b0ff7 /* 0x1ac8 */;
            1715: data_o = 32'h463341f7 /* 0x1acc */;
            1716: data_o = 32'he51700d7 /* 0x1ad0 */;
            1717: data_o = 32'he02effff /* 0x1ad4 */;
            1718: data_o = 32'h40d606bb /* 0x1ad8 */;
            1719: data_o = 32'h01f7571b /* 0x1adc */;
            1720: data_o = 32'h180c8626 /* 0x1ae0 */;
            1721: data_o = 32'h70e50513 /* 0x1ae4 */;
            1722: data_o = 32'hf693b755 /* 0x1ae8 */;
            1723: data_o = 32'hdef10806 /* 0x1aec */;
            1724: data_o = 32'h0107171b /* 0x1af0 */;
            1725: data_o = 32'h4107571b /* 0x1af4 */;
            1726: data_o = 32'hca99bfc9 /* 0x1af8 */;
            1727: data_o = 32'hffffe517 /* 0x1afc */;
            1728: data_o = 32'h47016014 /* 0x1b00 */;
            1729: data_o = 32'h8626e02e /* 0x1b04 */;
            1730: data_o = 32'h0513180c /* 0x1b08 */;
            1731: data_o = 32'hbfbd6e45 /* 0x1b0c */;
            1732: data_o = 32'h10077693 /* 0x1b10 */;
            1733: data_o = 32'he517ca99 /* 0x1b14 */;
            1734: data_o = 32'h6014ffff /* 0x1b18 */;
            1735: data_o = 32'he02e4701 /* 0x1b1c */;
            1736: data_o = 32'h180c8626 /* 0x1b20 */;
            1737: data_o = 32'h6ca50513 /* 0x1b24 */;
            1738: data_o = 32'h7613b795 /* 0x1b28 */;
            1739: data_o = 32'h40140407 /* 0x1b2c */;
            1740: data_o = 32'hf693ce11 /* 0x1b30 */;
            1741: data_o = 32'h16820ff6 /* 0x1b34 */;
            1742: data_o = 32'hffffe517 /* 0x1b38 */;
            1743: data_o = 32'h4701e02e /* 0x1b3c */;
            1744: data_o = 32'h86269281 /* 0x1b40 */;
            1745: data_o = 32'h0513180c /* 0x1b44 */;
            1746: data_o = 32'hb7896a85 /* 0x1b48 */;
            1747: data_o = 32'h08077713 /* 0x1b4c */;
            1748: data_o = 32'hf6b3d37d /* 0x1b50 */;
            1749: data_o = 32'hb7c50136 /* 0x1b54 */;
            1750: data_o = 32'h0205e593 /* 0x1b58 */;
            1751: data_o = 32'he5172008 /* 0x1b5c */;
            1752: data_o = 32'h87aeffff /* 0x1b60 */;
            1753: data_o = 32'h86c28746 /* 0x1b64 */;
            1754: data_o = 32'h180c8626 /* 0x1b68 */;
            1755: data_o = 32'h68250513 /* 0x1b6c */;
            1756: data_o = 32'h00840b93 /* 0x1b70 */;
            1757: data_o = 32'hbc0ff0ef /* 0x1b74 */;
            1758: data_o = 32'hfc13bf21 /* 0x1b78 */;
            1759: data_o = 32'h4b850025 /* 0x1b7c */;
            1760: data_o = 32'h040c1063 /* 0x1b80 */;
            1761: data_o = 32'ha8094b81 /* 0x1b84 */;
            1762: data_o = 32'h180c56fd /* 0x1b88 */;
            1763: data_o = 32'h02000513 /* 0x1b8c */;
            1764: data_o = 32'he0efec46 /* 0x1b90 */;
            1765: data_o = 32'h68e2e4ef /* 0x1b94 */;
            1766: data_o = 32'h01748633 /* 0x1b98 */;
            1767: data_o = 32'h879b0b85 /* 0x1b9c */;
            1768: data_o = 32'he3e3000b /* 0x1ba0 */;
            1769: data_o = 32'h4781ff17 /* 0x1ba4 */;
            1770: data_o = 32'h00088663 /* 0x1ba8 */;
            1771: data_o = 32'hfff8879b /* 0x1bac */;
            1772: data_o = 32'h93811782 /* 0x1bb0 */;
            1773: data_o = 32'h4b8994be /* 0x1bb4 */;
            1774: data_o = 32'h00088463 /* 0x1bb8 */;
            1775: data_o = 32'h00188b9b /* 0x1bbc */;
            1776: data_o = 32'h00044503 /* 0x1bc0 */;
            1777: data_o = 32'h862656fd /* 0x1bc4 */;
            1778: data_o = 32'hec46180c /* 0x1bc8 */;
            1779: data_o = 32'he14fe0ef /* 0x1bcc */;
            1780: data_o = 32'h0c9368e2 /* 0x1bd0 */;
            1781: data_o = 32'h8d130084 /* 0x1bd4 */;
            1782: data_o = 32'h0c630014 /* 0x1bd8 */;
            1783: data_o = 32'h845e020c /* 0x1bdc */;
            1784: data_o = 32'ha829866a /* 0x1be0 */;
            1785: data_o = 32'h180c56fd /* 0x1be4 */;
            1786: data_o = 32'h02000513 /* 0x1be8 */;
            1787: data_o = 32'h0493ec46 /* 0x1bec */;
            1788: data_o = 32'he0ef0016 /* 0x1bf0 */;
            1789: data_o = 32'h68e2deef /* 0x1bf4 */;
            1790: data_o = 32'h86262405 /* 0x1bf8 */;
            1791: data_o = 32'hff1464e3 /* 0x1bfc */;
            1792: data_o = 32'he7634781 /* 0x1c00 */;
            1793: data_o = 32'h8bbb0178 /* 0x1c04 */;
            1794: data_o = 32'h97934178 /* 0x1c08 */;
            1795: data_o = 32'h9381020b /* 0x1c0c */;
            1796: data_o = 32'h84669d3e /* 0x1c10 */;
            1797: data_o = 32'hbe0584ea /* 0x1c14 */;
            1798: data_o = 32'h00043d83 /* 0x1c18 */;
            1799: data_o = 32'h00840b93 /* 0x1c1c */;
            1800: data_o = 32'h056357fd /* 0x1c20 */;
            1801: data_o = 32'h17930008 /* 0x1c24 */;
            1802: data_o = 32'h93810208 /* 0x1c28 */;
            1803: data_o = 32'h8cee97ee /* 0x1c2c */;
            1804: data_o = 32'h0c85a011 /* 0x1c30 */;
            1805: data_o = 32'h000cc703 /* 0x1c34 */;
            1806: data_o = 32'h9ce3c319 /* 0x1c38 */;
            1807: data_o = 32'hfc13ff97 /* 0x1c3c */;
            1808: data_o = 32'h8cbb4005 /* 0x1c40 */;
            1809: data_o = 32'h086341bc /* 0x1c44 */;
            1810: data_o = 32'h87c2000c /* 0x1c48 */;
            1811: data_o = 32'h010cf363 /* 0x1c4c */;
            1812: data_o = 32'h8c9b87e6 /* 0x1c50 */;
            1813: data_o = 32'hf4130007 /* 0x1c54 */;
            1814: data_o = 32'he8210025 /* 0x1c58 */;
            1815: data_o = 32'h8d3b8626 /* 0x1c5c */;
            1816: data_o = 32'ha005409c /* 0x1c60 */;
            1817: data_o = 32'h00160793 /* 0x1c64 */;
            1818: data_o = 32'h180c56fd /* 0x1c68 */;
            1819: data_o = 32'h02000513 /* 0x1c6c */;
            1820: data_o = 32'hf042f446 /* 0x1c70 */;
            1821: data_o = 32'he0efec3e /* 0x1c74 */;
            1822: data_o = 32'h67e2d6af /* 0x1c78 */;
            1823: data_o = 32'h78a27802 /* 0x1c7c */;
            1824: data_o = 32'h07bb863e /* 0x1c80 */;
            1825: data_o = 32'hefe300cd /* 0x1c84 */;
            1826: data_o = 32'h873bfd17 /* 0x1c88 */;
            1827: data_o = 32'h47814198 /* 0x1c8c */;
            1828: data_o = 32'h0198e563 /* 0x1c90 */;
            1829: data_o = 32'h02071793 /* 0x1c94 */;
            1830: data_o = 32'h94be9381 /* 0x1c98 */;
            1831: data_o = 32'he3634781 /* 0x1c9c */;
            1832: data_o = 32'h87ba0198 /* 0x1ca0 */;
            1833: data_o = 32'h8cbb2c85 /* 0x1ca4 */;
            1834: data_o = 32'h8d260197 /* 0x1ca8 */;
            1835: data_o = 32'h883ea005 /* 0x1cac */;
            1836: data_o = 32'h001d0793 /* 0x1cb0 */;
            1837: data_o = 32'h56fd866a /* 0x1cb4 */;
            1838: data_o = 32'hf446180c /* 0x1cb8 */;
            1839: data_o = 32'hec3ef042 /* 0x1cbc */;
            1840: data_o = 32'hd20fe0ef /* 0x1cc0 */;
            1841: data_o = 32'h780267e2 /* 0x1cc4 */;
            1842: data_o = 32'h8d3e78a2 /* 0x1cc8 */;
            1843: data_o = 32'h409d07b3 /* 0x1ccc */;
            1844: data_o = 32'hc50397ee /* 0x1cd0 */;
            1845: data_o = 32'hc5190007 /* 0x1cd4 */;
            1846: data_o = 32'hfc0c0ce3 /* 0x1cd8 */;
            1847: data_o = 32'hfff8079b /* 0x1cdc */;
            1848: data_o = 32'hfc0817e3 /* 0x1ce0 */;
            1849: data_o = 32'h866acc0d /* 0x1ce4 */;
            1850: data_o = 32'h41ac843b /* 0x1ce8 */;
            1851: data_o = 32'h56fda821 /* 0x1cec */;
            1852: data_o = 32'h0513180c /* 0x1cf0 */;
            1853: data_o = 32'hec460200 /* 0x1cf4 */;
            1854: data_o = 32'h00160493 /* 0x1cf8 */;
            1855: data_o = 32'hce4fe0ef /* 0x1cfc */;
            1856: data_o = 32'h862668e2 /* 0x1d00 */;
            1857: data_o = 32'h00c407bb /* 0x1d04 */;
            1858: data_o = 32'hff17e3e3 /* 0x1d08 */;
            1859: data_o = 32'he7634781 /* 0x1d0c */;
            1860: data_o = 32'h8cbb0198 /* 0x1d10 */;
            1861: data_o = 32'h97934198 /* 0x1d14 */;
            1862: data_o = 32'h9381020c /* 0x1d18 */;
            1863: data_o = 32'h845e9d3e /* 0x1d1c */;
            1864: data_o = 32'h47a1bdd5 /* 0x1d20 */;
            1865: data_o = 32'h1101b311 /* 0x1d24 */;
            1866: data_o = 32'h0517e822 /* 0x1d28 */;
            1867: data_o = 32'he4170000 /* 0x1d2c */;
            1868: data_o = 32'h041300ff /* 0x1d30 */;
            1869: data_o = 32'h05132d24 /* 0x1d34 */;
            1870: data_o = 32'he42652e5 /* 0x1d38 */;
            1871: data_o = 32'hec06e04a /* 0x1d3c */;
            1872: data_o = 32'h00440913 /* 0x1d40 */;
            1873: data_o = 32'h9bdff0ef /* 0x1d44 */;
            1874: data_o = 32'h00840493 /* 0x1d48 */;
            1875: data_o = 32'h00042423 /* 0x1d4c */;
            1876: data_o = 32'hcf91409c /* 0x1d50 */;
            1877: data_o = 32'h00092783 /* 0x1d54 */;
            1878: data_o = 32'h100f2781 /* 0x1d58 */;
            1879: data_o = 32'h64420000 /* 0x1d5c */;
            1880: data_o = 32'h64a260e2 /* 0x1d60 */;
            1881: data_o = 32'h17826902 /* 0x1d64 */;
            1882: data_o = 32'h61059381 /* 0x1d68 */;
            1883: data_o = 32'h409c8782 /* 0x1d6c */;
            1884: data_o = 32'h0113b7c5 /* 0x1d70 */;
            1885: data_o = 32'h3823be01 /* 0x1d74 */;
            1886: data_o = 32'h34234081 /* 0x1d78 */;
            1887: data_o = 32'h30234091 /* 0x1d7c */;
            1888: data_o = 32'h84ae4121 /* 0x1d80 */;
            1889: data_o = 32'h4581842a /* 0x1d84 */;
            1890: data_o = 32'h00288932 /* 0x1d88 */;
            1891: data_o = 32'h1f800613 /* 0x1d8c */;
            1892: data_o = 32'h40113c23 /* 0x1d90 */;
            1893: data_o = 32'he0efe002 /* 0x1d94 */;
            1894: data_o = 32'h0613c24f /* 0x1d98 */;
            1895: data_o = 32'h45811f80 /* 0x1d9c */;
            1896: data_o = 32'h30230428 /* 0x1da0 */;
            1897: data_o = 32'he0ef2001 /* 0x1da4 */;
            1898: data_o = 32'h4685c14f /* 0x1da8 */;
            1899: data_o = 32'h4585860a /* 0x1dac */;
            1900: data_o = 32'h94028526 /* 0x1db0 */;
            1901: data_o = 32'h0517c115 /* 0x1db4 */;
            1902: data_o = 32'h05130000 /* 0x1db8 */;
            1903: data_o = 32'hf0ef4f25 /* 0x1dbc */;
            1904: data_o = 32'h3083943f /* 0x1dc0 */;
            1905: data_o = 32'h34034181 /* 0x1dc4 */;
            1906: data_o = 32'h34834101 /* 0x1dc8 */;
            1907: data_o = 32'h39034081 /* 0x1dcc */;
            1908: data_o = 32'h01134001 /* 0x1dd0 */;
            1909: data_o = 32'h80824201 /* 0x1dd4 */;
            1910: data_o = 32'h468545a6 /* 0x1dd8 */;
            1911: data_o = 32'h85260410 /* 0x1ddc */;
            1912: data_o = 32'hc5119402 /* 0x1de0 */;
            1913: data_o = 32'h00000517 /* 0x1de4 */;
            1914: data_o = 32'h4e450513 /* 0x1de8 */;
            1915: data_o = 32'h3783bfc9 /* 0x1dec */;
            1916: data_o = 32'h20232201 /* 0x1df0 */;
            1917: data_o = 32'hb7f100f9 /* 0x1df4 */;
            1918: data_o = 32'hf0a27159 /* 0x1df8 */;
            1919: data_o = 32'h00ffe417 /* 0x1dfc */;
            1920: data_o = 32'h20440413 /* 0x1e00 */;
            1921: data_o = 32'h27b75418 /* 0x1e04 */;
            1922: data_o = 32'hf486001c /* 0x1e08 */;
            1923: data_o = 32'h02f7573b /* 0x1e0c */;
            1924: data_o = 32'h01001797 /* 0x1e10 */;
            1925: data_o = 32'he8caeca6 /* 0x1e14 */;
            1926: data_o = 32'he0d2e4ce /* 0x1e18 */;
            1927: data_o = 32'h8793fc56 /* 0x1e1c */;
            1928: data_o = 32'h82231f07 /* 0x1e20 */;
            1929: data_o = 32'h06930007 /* 0x1e24 */;
            1930: data_o = 32'h8623f800 /* 0x1e28 */;
            1931: data_o = 32'h169700d7 /* 0x1e2c */;
            1932: data_o = 32'h76130100 /* 0x1e30 */;
            1933: data_o = 32'h571b0ff7 /* 0x1e34 */;
            1934: data_o = 32'h89230087 /* 0x1e38 */;
            1935: data_o = 32'h77131cc6 /* 0x1e3c */;
            1936: data_o = 32'h82230ff7 /* 0x1e40 */;
            1937: data_o = 32'h470d00e7 /* 0x1e44 */;
            1938: data_o = 32'h00e78623 /* 0x1e48 */;
            1939: data_o = 32'hfc700693 /* 0x1e4c */;
            1940: data_o = 32'h00d78423 /* 0x1e50 */;
            1941: data_o = 32'h02000693 /* 0x1e54 */;
            1942: data_o = 32'h00d78823 /* 0x1e58 */;
            1943: data_o = 32'h46894850 /* 0x1e5c */;
            1944: data_o = 32'h1ed60563 /* 0x1e60 */;
            1945: data_o = 32'h0006079b /* 0x1e64 */;
            1946: data_o = 32'h02840493 /* 0x1e68 */;
            1947: data_o = 32'h00f6ec63 /* 0x1e6c */;
            1948: data_o = 32'h0517e795 /* 0x1e70 */;
            1949: data_o = 32'h05130000 /* 0x1e74 */;
            1950: data_o = 32'hf0ef47e5 /* 0x1e78 */;
            1951: data_o = 32'hf0ef887f /* 0x1e7c */;
            1952: data_o = 32'ha2c9ea9f /* 0x1e80 */;
            1953: data_o = 32'h24e78163 /* 0x1e84 */;
            1954: data_o = 32'h01440593 /* 0x1e88 */;
            1955: data_o = 32'h0517418c /* 0x1e8c */;
            1956: data_o = 32'h05130000 /* 0x1e90 */;
            1957: data_o = 32'hf0ef52a5 /* 0x1e94 */;
            1958: data_o = 32'hb7d586bf /* 0x1e98 */;
            1959: data_o = 32'h00000517 /* 0x1e9c */;
            1960: data_o = 32'h47c50513 /* 0x1ea0 */;
            1961: data_o = 32'h85dff0ef /* 0x1ea4 */;
            1962: data_o = 32'h3717409c /* 0x1ea8 */;
            1963: data_o = 32'hec020100 /* 0x1eac */;
            1964: data_o = 32'h0007869b /* 0x1eb0 */;
            1965: data_o = 32'h15670713 /* 0x1eb4 */;
            1966: data_o = 32'hf402f002 /* 0x1eb8 */;
            1967: data_o = 32'he83ac202 /* 0x1ebc */;
            1968: data_o = 32'hd61bcc36 /* 0x1ec0 */;
            1969: data_o = 32'hd79b0017 /* 0x1ec4 */;
            1970: data_o = 32'hc2990017 /* 0x1ec8 */;
            1971: data_o = 32'hce32c3bd /* 0x1ecc */;
            1972: data_o = 32'hf0ef0808 /* 0x1ed0 */;
            1973: data_o = 32'h25b7b5ef /* 0x1ed4 */;
            1974: data_o = 32'h85930006 /* 0x1ed8 */;
            1975: data_o = 32'h0808a805 /* 0x1edc */;
            1976: data_o = 32'haf8ff0ef /* 0x1ee0 */;
            1977: data_o = 32'h04134985 /* 0x1ee4 */;
            1978: data_o = 32'h08080770 /* 0x1ee8 */;
            1979: data_o = 32'h02e99a13 /* 0x1eec */;
            1980: data_o = 32'h14225afd /* 0x1ef0 */;
            1981: data_o = 32'habaff0ef /* 0x1ef4 */;
            1982: data_o = 32'h0a134929 /* 0x1ef8 */;
            1983: data_o = 32'hda93095a /* 0x1efc */;
            1984: data_o = 32'h0413018a /* 0x1f00 */;
            1985: data_o = 32'h46010654 /* 0x1f04 */;
            1986: data_o = 32'h05000593 /* 0x1f08 */;
            1987: data_o = 32'he4020808 /* 0x1f0c */;
            1988: data_o = 32'haeefe0ef /* 0x1f10 */;
            1989: data_o = 32'h4681e149 /* 0x1f14 */;
            1990: data_o = 32'h85d20030 /* 0x1f18 */;
            1991: data_o = 32'hf0ef0808 /* 0x1f1c */;
            1992: data_o = 32'he935b66f /* 0x1f20 */;
            1993: data_o = 32'h00814783 /* 0x1f24 */;
            1994: data_o = 32'h01378b63 /* 0x1f28 */;
            1995: data_o = 32'he7a52781 /* 0x1f2c */;
            1996: data_o = 32'ha7b7a8d9 /* 0x1f30 */;
            1997: data_o = 32'h87930007 /* 0x1f34 */;
            1998: data_o = 32'hce3e1207 /* 0x1f38 */;
            1999: data_o = 32'h0797bf51 /* 0x1f3c */;
            2000: data_o = 32'hb5830000 /* 0x1f40 */;
            2001: data_o = 32'h469d5ea7 /* 0x1f44 */;
            2002: data_o = 32'h08080030 /* 0x1f48 */;
            2003: data_o = 32'hf0efe402 /* 0x1f4c */;
            2004: data_o = 32'he131b36f /* 0x1f50 */;
            2005: data_o = 32'h971367a2 /* 0x1f54 */;
            2006: data_o = 32'h07130209 /* 0x1f58 */;
            2007: data_o = 32'hf6b31aa7 /* 0x1f5c */;
            2008: data_o = 32'hf7930157 /* 0x1f60 */;
            2009: data_o = 32'h94e30ff7 /* 0x1f64 */;
            2010: data_o = 32'h4681fce6 /* 0x1f68 */;
            2011: data_o = 32'h85a20030 /* 0x1f6c */;
            2012: data_o = 32'he4020808 /* 0x1f70 */;
            2013: data_o = 32'hb10ff0ef /* 0x1f74 */;
            2014: data_o = 32'h0493ed19 /* 0x1f78 */;
            2015: data_o = 32'h149a1a50 /* 0x1f7c */;
            2016: data_o = 32'h07748593 /* 0x1f80 */;
            2017: data_o = 32'h00304681 /* 0x1f84 */;
            2018: data_o = 32'he4020808 /* 0x1f88 */;
            2019: data_o = 32'haf8ff0ef /* 0x1f8c */;
            2020: data_o = 32'h07748493 /* 0x1f90 */;
            2021: data_o = 32'h397dcd05 /* 0x1f94 */;
            2022: data_o = 32'hf60917e3 /* 0x1f98 */;
            2023: data_o = 32'h00000517 /* 0x1f9c */;
            2024: data_o = 32'h45c50513 /* 0x1fa0 */;
            2025: data_o = 32'hf5cff0ef /* 0x1fa4 */;
            2026: data_o = 32'hd7fff0ef /* 0x1fa8 */;
            2027: data_o = 32'h4681a8a9 /* 0x1fac */;
            2028: data_o = 32'h85a20030 /* 0x1fb0 */;
            2029: data_o = 32'hf0ef0808 /* 0x1fb4 */;
            2030: data_o = 32'hfd71acef /* 0x1fb8 */;
            2031: data_o = 32'h00304681 /* 0x1fbc */;
            2032: data_o = 32'h080885a6 /* 0x1fc0 */;
            2033: data_o = 32'hf0efe402 /* 0x1fc4 */;
            2034: data_o = 32'hf571abef /* 0x1fc8 */;
            2035: data_o = 32'h00814783 /* 0x1fcc */;
            2036: data_o = 32'hfff1e402 /* 0x1fd0 */;
            2037: data_o = 32'h03d00593 /* 0x1fd4 */;
            2038: data_o = 32'h468d15a6 /* 0x1fd8 */;
            2039: data_o = 32'h85930030 /* 0x1fdc */;
            2040: data_o = 32'h08080fd5 /* 0x1fe0 */;
            2041: data_o = 32'haa0ff0ef /* 0x1fe4 */;
            2042: data_o = 32'h0797f55d /* 0x1fe8 */;
            2043: data_o = 32'hb5830000 /* 0x1fec */;
            2044: data_o = 32'h46815467 /* 0x1ff0 */;
            2045: data_o = 32'h08080030 /* 0x1ff4 */;
            2046: data_o = 32'hf0efe402 /* 0x1ff8 */;
            2047: data_o = 32'hfd41a8af /* 0x1ffc */;
            2048: data_o = 32'h00814783 /* 0x2000 */;
            2049: data_o = 32'hc5b7f785 /* 0x2004 */;
            2050: data_o = 32'h859300be /* 0x2008 */;
            2051: data_o = 32'h0808c205 /* 0x200c */;
            2052: data_o = 32'h9c8ff0ef /* 0x2010 */;
            2053: data_o = 32'hfffff517 /* 0x2014 */;
            2054: data_o = 32'h080c0050 /* 0x2018 */;
            2055: data_o = 32'h6e450513 /* 0x201c */;
            2056: data_o = 32'hd53ff0ef /* 0x2020 */;
            2057: data_o = 32'he6174592 /* 0x2024 */;
            2058: data_o = 32'h06936eff /* 0x2028 */;
            2059: data_o = 32'h06130200 /* 0x202c */;
            2060: data_o = 32'h0808fda6 /* 0x2030 */;
            2061: data_o = 32'hba8ff0ef /* 0x2034 */;
            2062: data_o = 32'h0000100f /* 0x2038 */;
            2063: data_o = 32'h6effe097 /* 0x203c */;
            2064: data_o = 32'hfc4080e7 /* 0x2040 */;
            2065: data_o = 32'h10500073 /* 0x2044 */;
            2066: data_o = 32'h0517bff5 /* 0x2048 */;
            2067: data_o = 32'h05130000 /* 0x204c */;
            2068: data_o = 32'hf0ef2fe5 /* 0x2050 */;
            2069: data_o = 32'h541ceaef /* 0x2054 */;
            2070: data_o = 32'h01003717 /* 0x2058 */;
            2071: data_o = 32'h869bec02 /* 0x205c */;
            2072: data_o = 32'h07130007 /* 0x2060 */;
            2073: data_o = 32'hf002fa87 /* 0x2064 */;
            2074: data_o = 32'hc402f402 /* 0x2068 */;
            2075: data_o = 32'hcc36e83a /* 0x206c */;
            2076: data_o = 32'h0017d79b /* 0x2070 */;
            2077: data_o = 32'he789ca89 /* 0x2074 */;
            2078: data_o = 32'h0007a7b7 /* 0x2078 */;
            2079: data_o = 32'h12078793 /* 0x207c */;
            2080: data_o = 32'h4785ce3e /* 0x2080 */;
            2081: data_o = 32'h0808d03e /* 0x2084 */;
            2082: data_o = 32'h9a8ff0ef /* 0x2088 */;
            2083: data_o = 32'h017d85b7 /* 0x208c */;
            2084: data_o = 32'h84058593 /* 0x2090 */;
            2085: data_o = 32'hf0ef0808 /* 0x2094 */;
            2086: data_o = 32'h0808942f /* 0x2098 */;
            2087: data_o = 32'h912ff0ef /* 0x209c */;
            2088: data_o = 32'hffffe517 /* 0x20a0 */;
            2089: data_o = 32'h080c0030 /* 0x20a4 */;
            2090: data_o = 32'h6d050513 /* 0x20a8 */;
            2091: data_o = 32'hcc7ff0ef /* 0x20ac */;
            2092: data_o = 32'he61745a2 /* 0x20b0 */;
            2093: data_o = 32'h06936eff /* 0x20b4 */;
            2094: data_o = 32'h06130200 /* 0x20b8 */;
            2095: data_o = 32'h0808f4e6 /* 0x20bc */;
            2096: data_o = 32'he36fe0ef /* 0x20c0 */;
            2097: data_o = 32'h0517bf95 /* 0x20c4 */;
            2098: data_o = 32'h05130000 /* 0x20c8 */;
            2099: data_o = 32'hf0ef2b25 /* 0x20cc */;
            2100: data_o = 32'h409ce32f /* 0x20d0 */;
            2101: data_o = 32'h3b9ad537 /* 0x20d4 */;
            2102: data_o = 32'ha005051b /* 0x20d8 */;
            2103: data_o = 32'h02f5553b /* 0x20dc */;
            2104: data_o = 32'h3e700693 /* 0x20e0 */;
            2105: data_o = 32'h12b00613 /* 0x20e4 */;
            2106: data_o = 32'h05936705 /* 0x20e8 */;
            2107: data_o = 32'h071b5130 /* 0x20ec */;
            2108: data_o = 32'h2797bba7 /* 0x20f0 */;
            2109: data_o = 32'h87930100 /* 0x20f4 */;
            2110: data_o = 32'he83ef0e7 /* 0x20f8 */;
            2111: data_o = 32'h25700793 /* 0x20fc */;
            2112: data_o = 32'hd6bbc402 /* 0x2100 */;
            2113: data_o = 32'h563b02a6 /* 0x2104 */;
            2114: data_o = 32'h268502a6 /* 0x2108 */;
            2115: data_o = 32'h92c116c2 /* 0x210c */;
            2116: data_o = 32'h02a5d5bb /* 0x2110 */;
            2117: data_o = 32'h16422605 /* 0x2114 */;
            2118: data_o = 32'h573b9241 /* 0x2118 */;
            2119: data_o = 32'h881b02a7 /* 0x211c */;
            2120: data_o = 32'h181b0015 /* 0x2120 */;
            2121: data_o = 32'hd7bb0108 /* 0x2124 */;
            2122: data_o = 32'h9f0d02a7 /* 0x2128 */;
            2123: data_o = 32'h9f119f15 /* 0x212c */;
            2124: data_o = 32'h174285ba /* 0x2130 */;
            2125: data_o = 32'h27859341 /* 0x2134 */;
            2126: data_o = 32'h03079893 /* 0x2138 */;
            2127: data_o = 32'h7ff7f793 /* 0x213c */;
            2128: data_o = 32'h0308d893 /* 0x2140 */;
            2129: data_o = 32'h00f77363 /* 0x2144 */;
            2130: data_o = 32'h959b85c6 /* 0x2148 */;
            2131: data_o = 32'hd59b0105 /* 0x214c */;
            2132: data_o = 32'he5b30105 /* 0x2150 */;
            2133: data_o = 32'h27170105 /* 0x2154 */;
            2134: data_o = 32'h25810100 /* 0x2158 */;
            2135: data_o = 32'heaa70713 /* 0x215c */;
            2136: data_o = 32'h0106161b /* 0x2160 */;
            2137: data_o = 32'h8ed1db0c /* 0x2164 */;
            2138: data_o = 32'h01002717 /* 0x2168 */;
            2139: data_o = 32'h07132681 /* 0x216c */;
            2140: data_o = 32'hdb54e987 /* 0x2170 */;
            2141: data_o = 32'h01079693 /* 0x2174 */;
            2142: data_o = 32'h01002717 /* 0x2178 */;
            2143: data_o = 32'h07138edd /* 0x217c */;
            2144: data_o = 32'hdf14e887 /* 0x2180 */;
            2145: data_o = 32'h06300713 /* 0x2184 */;
            2146: data_o = 32'h02a7573b /* 0x2188 */;
            2147: data_o = 32'he7b366c1 /* 0x218c */;
            2148: data_o = 32'h27810107 /* 0x2190 */;
            2149: data_o = 32'h45814605 /* 0x2194 */;
            2150: data_o = 32'h8f552705 /* 0x2198 */;
            2151: data_o = 32'h01002697 /* 0x219c */;
            2152: data_o = 32'he6468693 /* 0x21a0 */;
            2153: data_o = 32'hded82701 /* 0x21a4 */;
            2154: data_o = 32'h01002717 /* 0x21a8 */;
            2155: data_o = 32'he5870713 /* 0x21ac */;
            2156: data_o = 32'h2797c33c /* 0x21b0 */;
            2157: data_o = 32'h87930100 /* 0x21b4 */;
            2158: data_o = 32'h4b88e4e7 /* 0x21b8 */;
            2159: data_o = 32'hdb6fe0ef /* 0x21bc */;
            2160: data_o = 32'h01002797 /* 0x21c0 */;
            2161: data_o = 32'he4078793 /* 0x21c4 */;
            2162: data_o = 32'hcb882501 /* 0x21c8 */;
            2163: data_o = 32'hfffff517 /* 0x21cc */;
            2164: data_o = 32'h080c0030 /* 0x21d0 */;
            2165: data_o = 32'h82450513 /* 0x21d4 */;
            2166: data_o = 32'hb9bff0ef /* 0x21d8 */;
            2167: data_o = 32'he61745a2 /* 0x21dc */;
            2168: data_o = 32'h06936eff /* 0x21e0 */;
            2169: data_o = 32'h06130200 /* 0x21e4 */;
            2170: data_o = 32'h0808e226 /* 0x21e8 */;
            2171: data_o = 32'he3efe0ef /* 0x21ec */;
            2172: data_o = 32'h0000b5a1 /* 0x21f0 */;
            2173: data_o = 32'h00000000 /* 0x21f4 */;
            2174: data_o = 32'h2b696e66 /* 0x21f8 */;
            2175: data_o = 32'h00000000 /* 0x21fc */;
            2176: data_o = 32'h00696e66 /* 0x2200 */;
            2177: data_o = 32'h00000000 /* 0x2204 */;
            2178: data_o = 32'h006e616e /* 0x2208 */;
            2179: data_o = 32'h00000000 /* 0x220c */;
            2180: data_o = 32'h2d696e66 /* 0x2210 */;
            2181: data_o = 32'h00000000 /* 0x2214 */;
            2182: data_o = 32'hfffff7f4 /* 0x2218 */;
            2183: data_o = 32'hfffff570 /* 0x221c */;
            2184: data_o = 32'hfffff570 /* 0x2220 */;
            2185: data_o = 32'hfffff570 /* 0x2224 */;
            2186: data_o = 32'hfffff570 /* 0x2228 */;
            2187: data_o = 32'hfffff570 /* 0x222c */;
            2188: data_o = 32'hfffff570 /* 0x2230 */;
            2189: data_o = 32'hfffff570 /* 0x2234 */;
            2190: data_o = 32'hfffff570 /* 0x2238 */;
            2191: data_o = 32'hfffff570 /* 0x223c */;
            2192: data_o = 32'hfffff7f4 /* 0x2240 */;
            2193: data_o = 32'hfffff962 /* 0x2244 */;
            2194: data_o = 32'hfffff7f4 /* 0x2248 */;
            2195: data_o = 32'hfffff766 /* 0x224c */;
            2196: data_o = 32'hfffff944 /* 0x2250 */;
            2197: data_o = 32'hfffff766 /* 0x2254 */;
            2198: data_o = 32'h6f6f625b /* 0x2258 */;
            2199: data_o = 32'h6d6f7274 /* 0x225c */;
            2200: data_o = 32'h6f50205d /* 0x2260 */;
            2201: data_o = 32'h6e696c6c /* 0x2264 */;
            2202: data_o = 32'h63732067 /* 0x2268 */;
            2203: data_o = 32'h63746172 /* 0x226c */;
            2204: data_o = 32'h66203068 /* 0x2270 */;
            2205: data_o = 32'h6520726f /* 0x2274 */;
            2206: data_o = 32'h7972746e /* 0x2278 */;
            2207: data_o = 32'h696f7020 /* 0x227c */;
            2208: data_o = 32'h6120746e /* 0x2280 */;
            2209: data_o = 32'h7320646e /* 0x2284 */;
            2210: data_o = 32'h74617263 /* 0x2288 */;
            2211: data_o = 32'h20316863 /* 0x228c */;
            2212: data_o = 32'h20726f66 /* 0x2290 */;
            2213: data_o = 32'h72617473 /* 0x2294 */;
            2214: data_o = 32'h69732074 /* 0x2298 */;
            2215: data_o = 32'h6c616e67 /* 0x229c */;
            2216: data_o = 32'h000a0d2e /* 0x22a0 */;
            2217: data_o = 32'h00000000 /* 0x22a4 */;
            2218: data_o = 32'h79706f43 /* 0x22a8 */;
            2219: data_o = 32'h20676e69 /* 0x22ac */;
            2220: data_o = 32'h20656874 /* 0x22b0 */;
            2221: data_o = 32'h64616568 /* 0x22b4 */;
            2222: data_o = 32'h66207265 /* 0x22b8 */;
            2223: data_o = 32'h656c6961 /* 0x22bc */;
            2224: data_o = 32'h0a0d2164 /* 0x22c0 */;
            2225: data_o = 32'h00000000 /* 0x22c4 */;
            2226: data_o = 32'h79706f43 /* 0x22c8 */;
            2227: data_o = 32'h20676e69 /* 0x22cc */;
            2228: data_o = 32'h20656874 /* 0x22d0 */;
            2229: data_o = 32'h74726170 /* 0x22d4 */;
            2230: data_o = 32'h6f697469 /* 0x22d8 */;
            2231: data_o = 32'h6e65206e /* 0x22dc */;
            2232: data_o = 32'h65697274 /* 0x22e0 */;
            2233: data_o = 32'h61662073 /* 0x22e4 */;
            2234: data_o = 32'h64656c69 /* 0x22e8 */;
            2235: data_o = 32'h000a0d21 /* 0x22ec */;
            2236: data_o = 32'h6f6f625b /* 0x22f0 */;
            2237: data_o = 32'h6d6f7274 /* 0x22f4 */;
            2238: data_o = 32'h6f42205d /* 0x22f8 */;
            2239: data_o = 32'h6f6d746f /* 0x22fc */;
            2240: data_o = 32'h30206564 /* 0x2300 */;
            2241: data_o = 32'h6449203a /* 0x2304 */;
            2242: data_o = 32'h6220656c /* 0x2308 */;
            2243: data_o = 32'h2e746f6f /* 0x230c */;
            2244: data_o = 32'h00000a0d /* 0x2310 */;
            2245: data_o = 32'h00000000 /* 0x2314 */;
            2246: data_o = 32'h6f6f625b /* 0x2318 */;
            2247: data_o = 32'h6d6f7274 /* 0x231c */;
            2248: data_o = 32'h6f42205d /* 0x2320 */;
            2249: data_o = 32'h6f6d746f /* 0x2324 */;
            2250: data_o = 32'h31206564 /* 0x2328 */;
            2251: data_o = 32'h4453203a /* 0x232c */;
            2252: data_o = 32'h72616320 /* 0x2330 */;
            2253: data_o = 32'h6f622064 /* 0x2334 */;
            2254: data_o = 32'h2820746f /* 0x2338 */;
            2255: data_o = 32'h30205343 /* 0x233c */;
            2256: data_o = 32'h000a0d29 /* 0x2340 */;
            2257: data_o = 32'h00000000 /* 0x2344 */;
            2258: data_o = 32'h6f6f625b /* 0x2348 */;
            2259: data_o = 32'h6d6f7274 /* 0x234c */;
            2260: data_o = 32'h6f42205d /* 0x2350 */;
            2261: data_o = 32'h6f6d746f /* 0x2354 */;
            2262: data_o = 32'h32206564 /* 0x2358 */;
            2263: data_o = 32'h5053203a /* 0x235c */;
            2264: data_o = 32'h6c662049 /* 0x2360 */;
            2265: data_o = 32'h20687361 /* 0x2364 */;
            2266: data_o = 32'h746f6f62 /* 0x2368 */;
            2267: data_o = 32'h53432820 /* 0x236c */;
            2268: data_o = 32'h0d293120 /* 0x2370 */;
            2269: data_o = 32'h0000000a /* 0x2374 */;
            2270: data_o = 32'h6f6f625b /* 0x2378 */;
            2271: data_o = 32'h6d6f7274 /* 0x237c */;
            2272: data_o = 32'h6f42205d /* 0x2380 */;
            2273: data_o = 32'h6f6d746f /* 0x2384 */;
            2274: data_o = 32'h33206564 /* 0x2388 */;
            2275: data_o = 32'h3249203a /* 0x238c */;
            2276: data_o = 32'h6c662043 /* 0x2390 */;
            2277: data_o = 32'h20687361 /* 0x2394 */;
            2278: data_o = 32'h746f6f62 /* 0x2398 */;
            2279: data_o = 32'h64612820 /* 0x239c */;
            2280: data_o = 32'h203a7264 /* 0x23a0 */;
            2281: data_o = 32'h30316230 /* 0x23a4 */;
            2282: data_o = 32'h30303031 /* 0x23a8 */;
            2283: data_o = 32'h0a0d2930 /* 0x23ac */;
            2284: data_o = 32'h00000000 /* 0x23b0 */;
            2285: data_o = 32'h00000000 /* 0x23b4 */;
            2286: data_o = 32'h6f6f625b /* 0x23b8 */;
            2287: data_o = 32'h6d6f7274 /* 0x23bc */;
            2288: data_o = 32'h6f42205d /* 0x23c0 */;
            2289: data_o = 32'h6f6d746f /* 0x23c4 */;
            2290: data_o = 32'h25206564 /* 0x23c8 */;
            2291: data_o = 32'h55203a64 /* 0x23cc */;
            2292: data_o = 32'h6f6e6b6e /* 0x23d0 */;
            2293: data_o = 32'h62206e77 /* 0x23d4 */;
            2294: data_o = 32'h6d746f6f /* 0x23d8 */;
            2295: data_o = 32'h2e65646f /* 0x23dc */;
            2296: data_o = 32'h69735520 /* 0x23e0 */;
            2297: data_o = 32'h6920676e /* 0x23e4 */;
            2298: data_o = 32'h20656c64 /* 0x23e8 */;
            2299: data_o = 32'h746f6f62 /* 0x23ec */;
            2300: data_o = 32'h000a0d2e /* 0x23f0 */;
            2301: data_o = 32'h00000000 /* 0x23f4 */;
            2302: data_o = 32'h6f6f625b /* 0x23f8 */;
            2303: data_o = 32'h6d6f7274 /* 0x23fc */;
            2304: data_o = 32'h6f43205d /* 0x2400 */;
            2305: data_o = 32'h20646c75 /* 0x2404 */;
            2306: data_o = 32'h20746f6e /* 0x2408 */;
            2307: data_o = 32'h74696e69 /* 0x240c */;
            2308: data_o = 32'h696c6169 /* 0x2410 */;
            2309: data_o = 32'h6120657a /* 0x2414 */;
            2310: data_o = 32'h20445320 /* 0x2418 */;
            2311: data_o = 32'h64726163 /* 0x241c */;
            2312: data_o = 32'h6146202e /* 0x2420 */;
            2313: data_o = 32'h6e696c6c /* 0x2424 */;
            2314: data_o = 32'h61622067 /* 0x2428 */;
            2315: data_o = 32'h74206b63 /* 0x242c */;
            2316: data_o = 32'h6469206f /* 0x2430 */;
            2317: data_o = 32'h6220656c /* 0x2434 */;
            2318: data_o = 32'h21746f6f /* 0x2438 */;
            2319: data_o = 32'h00000a0d /* 0x243c */;
            2320: data_o = 32'h00000000 /* 0x2440 */;
            2321: data_o = 32'h3ff00000 /* 0x2444 */;
            2322: data_o = 32'h00000000 /* 0x2448 */;
            2323: data_o = 32'h40240000 /* 0x244c */;
            2324: data_o = 32'h00000000 /* 0x2450 */;
            2325: data_o = 32'h40590000 /* 0x2454 */;
            2326: data_o = 32'h00000000 /* 0x2458 */;
            2327: data_o = 32'h408f4000 /* 0x245c */;
            2328: data_o = 32'h00000000 /* 0x2460 */;
            2329: data_o = 32'h40c38800 /* 0x2464 */;
            2330: data_o = 32'h00000000 /* 0x2468 */;
            2331: data_o = 32'h40f86a00 /* 0x246c */;
            2332: data_o = 32'h00000000 /* 0x2470 */;
            2333: data_o = 32'h412e8480 /* 0x2474 */;
            2334: data_o = 32'h00000000 /* 0x2478 */;
            2335: data_o = 32'h416312d0 /* 0x247c */;
            2336: data_o = 32'h00000000 /* 0x2480 */;
            2337: data_o = 32'h4197d784 /* 0x2484 */;
            2338: data_o = 32'h00000000 /* 0x2488 */;
            2339: data_o = 32'h41cdcd65 /* 0x248c */;
            2340: data_o = 32'hffffffff /* 0x2490 */;
            2341: data_o = 32'h7fefffff /* 0x2494 */;
            2342: data_o = 32'hffffffff /* 0x2498 */;
            2343: data_o = 32'hffefffff /* 0x249c */;
            2344: data_o = 32'h509f79fb /* 0x24a0 */;
            2345: data_o = 32'h3fd34413 /* 0x24a4 */;
            2346: data_o = 32'h8b60c8b3 /* 0x24a8 */;
            2347: data_o = 32'h3fc68a28 /* 0x24ac */;
            2348: data_o = 32'h00000000 /* 0x24b0 */;
            2349: data_o = 32'h3ff80000 /* 0x24b4 */;
            2350: data_o = 32'h636f4361 /* 0x24b8 */;
            2351: data_o = 32'h3fd287a7 /* 0x24bc */;
            2352: data_o = 32'h0979a371 /* 0x24c0 */;
            2353: data_o = 32'h400a934f /* 0x24c4 */;
            2354: data_o = 32'h00000000 /* 0x24c8 */;
            2355: data_o = 32'h3fe00000 /* 0x24cc */;
            2356: data_o = 32'hfefa39ef /* 0x24d0 */;
            2357: data_o = 32'h3fe62e42 /* 0x24d4 */;
            2358: data_o = 32'hbbb55516 /* 0x24d8 */;
            2359: data_o = 32'h40026bb1 /* 0x24dc */;
            2360: data_o = 32'h00000000 /* 0x24e0 */;
            2361: data_o = 32'h402c0000 /* 0x24e4 */;
            2362: data_o = 32'h00000000 /* 0x24e8 */;
            2363: data_o = 32'h40240000 /* 0x24ec */;
            2364: data_o = 32'h00000000 /* 0x24f0 */;
            2365: data_o = 32'h40180000 /* 0x24f4 */;
            2366: data_o = 32'h00000000 /* 0x24f8 */;
            2367: data_o = 32'h40000000 /* 0x24fc */;
            2368: data_o = 32'h00000000 /* 0x2500 */;
            2369: data_o = 32'h3ff00000 /* 0x2504 */;
            2370: data_o = 32'heb1c432d /* 0x2508 */;
            2371: data_o = 32'h3f1a36e2 /* 0x250c */;
            2372: data_o = 32'h00000000 /* 0x2510 */;
            2373: data_o = 32'h412e8480 /* 0x2514 */;
            2374: data_o = 32'h00000000 /* 0x2518 */;
            2375: data_o = 32'h41cdcd65 /* 0x251c */;
            2376: data_o = 32'h00000000 /* 0x2520 */;
            2377: data_o = 32'hc1cdcd65 /* 0x2524 */;
            2378: data_o = 32'h0001aa87 /* 0x2528 */;
            2379: data_o = 32'h00004800 /* 0x252c */;
            2380: data_o = 32'h00020015 /* 0x2530 */;
            2381: data_o = 32'h00005000 /* 0x2534 */;
            2382: data_o = 32'h05020101 /* 0x2538 */;
            2383: data_o = 32'h05000000 /* 0x253c */;
            2384: data_o = 32'h00000000 /* 0x2540 */;
            2385: data_o = 32'h00000000 /* 0x2544 */;
            2386: data_o = 32'h00000000 /* 0x2548 */;
            2387: data_o = 32'h00000000 /* 0x254c */;
            2388: data_o = 32'h00000000 /* 0x2550 */;
            2389: data_o = 32'h00000000 /* 0x2554 */;
            2390: data_o = 32'h00000000 /* 0x2558 */;
            2391: data_o = 32'h00000000 /* 0x255c */;
            2392: data_o = 32'h00000000 /* 0x2560 */;
            2393: data_o = 32'h00000000 /* 0x2564 */;
            2394: data_o = 32'h00000000 /* 0x2568 */;
            2395: data_o = 32'h00000000 /* 0x256c */;
            2396: data_o = 32'h00000000 /* 0x2570 */;
            2397: data_o = 32'h00000000 /* 0x2574 */;
            2398: data_o = 32'h00000000 /* 0x2578 */;
            2399: data_o = 32'h00000000 /* 0x257c */;
            2400: data_o = 32'h00000000 /* 0x2580 */;
            2401: data_o = 32'h00000000 /* 0x2584 */;
            2402: data_o = 32'h00000000 /* 0x2588 */;
            2403: data_o = 32'h00000000 /* 0x258c */;
            2404: data_o = 32'h00000000 /* 0x2590 */;
            2405: data_o = 32'h00000000 /* 0x2594 */;
            2406: data_o = 32'h00000000 /* 0x2598 */;
            2407: data_o = 32'h00000000 /* 0x259c */;
            2408: data_o = 32'h00000000 /* 0x25a0 */;
            2409: data_o = 32'h00000000 /* 0x25a4 */;
            2410: data_o = 32'h00000000 /* 0x25a8 */;
            2411: data_o = 32'h00000000 /* 0x25ac */;
            2412: data_o = 32'h00000000 /* 0x25b0 */;
            2413: data_o = 32'h00000000 /* 0x25b4 */;
            2414: data_o = 32'h00000000 /* 0x25b8 */;
            2415: data_o = 32'h00000000 /* 0x25bc */;
            2416: data_o = 32'h00000000 /* 0x25c0 */;
            2417: data_o = 32'h00000000 /* 0x25c4 */;
            2418: data_o = 32'h00000000 /* 0x25c8 */;
            2419: data_o = 32'h00000000 /* 0x25cc */;
            2420: data_o = 32'h00000000 /* 0x25d0 */;
            2421: data_o = 32'h00000000 /* 0x25d4 */;
            2422: data_o = 32'h00000000 /* 0x25d8 */;
            2423: data_o = 32'h00000000 /* 0x25dc */;
            2424: data_o = 32'h00000000 /* 0x25e0 */;
            2425: data_o = 32'h00000000 /* 0x25e4 */;
            2426: data_o = 32'h00000000 /* 0x25e8 */;
            2427: data_o = 32'h00000000 /* 0x25ec */;
            2428: data_o = 32'h00000000 /* 0x25f0 */;
            2429: data_o = 32'h00000000 /* 0x25f4 */;
            2430: data_o = 32'h00000000 /* 0x25f8 */;
            2431: data_o = 32'h00000000 /* 0x25fc */;
            2432: data_o = 32'h00000000 /* 0x2600 */;
            2433: data_o = 32'h00000000 /* 0x2604 */;
            2434: data_o = 32'h00000000 /* 0x2608 */;
            2435: data_o = 32'h00000000 /* 0x260c */;
            2436: data_o = 32'h00000000 /* 0x2610 */;
            2437: data_o = 32'h00000000 /* 0x2614 */;
            2438: data_o = 32'h00000000 /* 0x2618 */;
            2439: data_o = 32'h00000000 /* 0x261c */;
            2440: data_o = 32'h00000000 /* 0x2620 */;
            2441: data_o = 32'h00000000 /* 0x2624 */;
            2442: data_o = 32'h00000000 /* 0x2628 */;
            2443: data_o = 32'h00000000 /* 0x262c */;
            2444: data_o = 32'h00000000 /* 0x2630 */;
            2445: data_o = 32'h00000000 /* 0x2634 */;
            2446: data_o = 32'h00000000 /* 0x2638 */;
            2447: data_o = 32'h00000000 /* 0x263c */;
            2448: data_o = 32'h00000000 /* 0x2640 */;
            2449: data_o = 32'h00000000 /* 0x2644 */;
            2450: data_o = 32'h00000000 /* 0x2648 */;
            2451: data_o = 32'h00000000 /* 0x264c */;
            2452: data_o = 32'h00000000 /* 0x2650 */;
            2453: data_o = 32'h00000000 /* 0x2654 */;
            2454: data_o = 32'h00000000 /* 0x2658 */;
            2455: data_o = 32'h00000000 /* 0x265c */;
            2456: data_o = 32'h00000000 /* 0x2660 */;
            2457: data_o = 32'h00000000 /* 0x2664 */;
            2458: data_o = 32'h00000000 /* 0x2668 */;
            2459: data_o = 32'h00000000 /* 0x266c */;
            2460: data_o = 32'h00000000 /* 0x2670 */;
            2461: data_o = 32'h00000000 /* 0x2674 */;
            2462: data_o = 32'h00000000 /* 0x2678 */;
            2463: data_o = 32'h00000000 /* 0x267c */;
            2464: data_o = 32'h00000000 /* 0x2680 */;
            2465: data_o = 32'h00000000 /* 0x2684 */;
            2466: data_o = 32'h00000000 /* 0x2688 */;
            2467: data_o = 32'h00000000 /* 0x268c */;
            2468: data_o = 32'h00000000 /* 0x2690 */;
            2469: data_o = 32'h00000000 /* 0x2694 */;
            2470: data_o = 32'h00000000 /* 0x2698 */;
            2471: data_o = 32'h00000000 /* 0x269c */;
            2472: data_o = 32'h00000000 /* 0x26a0 */;
            2473: data_o = 32'h00000000 /* 0x26a4 */;
            2474: data_o = 32'h00000000 /* 0x26a8 */;
            2475: data_o = 32'h00000000 /* 0x26ac */;
            2476: data_o = 32'h00000000 /* 0x26b0 */;
            2477: data_o = 32'h00000000 /* 0x26b4 */;
            2478: data_o = 32'h00000000 /* 0x26b8 */;
            2479: data_o = 32'h00000000 /* 0x26bc */;
            2480: data_o = 32'h00000000 /* 0x26c0 */;
            2481: data_o = 32'h00000000 /* 0x26c4 */;
            2482: data_o = 32'h00000000 /* 0x26c8 */;
            2483: data_o = 32'h00000000 /* 0x26cc */;
            2484: data_o = 32'h00000000 /* 0x26d0 */;
            2485: data_o = 32'h00000000 /* 0x26d4 */;
            2486: data_o = 32'h00000000 /* 0x26d8 */;
            2487: data_o = 32'h00000000 /* 0x26dc */;
            2488: data_o = 32'h00000000 /* 0x26e0 */;
            2489: data_o = 32'h00000000 /* 0x26e4 */;
            2490: data_o = 32'h00000000 /* 0x26e8 */;
            2491: data_o = 32'h00000000 /* 0x26ec */;
            2492: data_o = 32'h00000000 /* 0x26f0 */;
            2493: data_o = 32'h00000000 /* 0x26f4 */;
            2494: data_o = 32'h00000000 /* 0x26f8 */;
            2495: data_o = 32'h00000000 /* 0x26fc */;
            2496: data_o = 32'h00000000 /* 0x2700 */;
            2497: data_o = 32'h00000000 /* 0x2704 */;
            2498: data_o = 32'h00000000 /* 0x2708 */;
            2499: data_o = 32'h00000000 /* 0x270c */;
            2500: data_o = 32'h00000000 /* 0x2710 */;
            2501: data_o = 32'h00000000 /* 0x2714 */;
            2502: data_o = 32'h00000000 /* 0x2718 */;
            2503: data_o = 32'h00000000 /* 0x271c */;
            2504: data_o = 32'h00000000 /* 0x2720 */;
            2505: data_o = 32'h00000000 /* 0x2724 */;
            2506: data_o = 32'h00000000 /* 0x2728 */;
            2507: data_o = 32'h00000000 /* 0x272c */;
            2508: data_o = 32'h00000000 /* 0x2730 */;
            2509: data_o = 32'h00000000 /* 0x2734 */;
            2510: data_o = 32'h00000000 /* 0x2738 */;
            2511: data_o = 32'h00000000 /* 0x273c */;
            2512: data_o = 32'h00000000 /* 0x2740 */;
            2513: data_o = 32'h00000000 /* 0x2744 */;
            2514: data_o = 32'h00000000 /* 0x2748 */;
            2515: data_o = 32'h00000000 /* 0x274c */;
            2516: data_o = 32'h00000000 /* 0x2750 */;
            2517: data_o = 32'h00000000 /* 0x2754 */;
            2518: data_o = 32'h00000000 /* 0x2758 */;
            2519: data_o = 32'h00000000 /* 0x275c */;
            2520: data_o = 32'h00000000 /* 0x2760 */;
            2521: data_o = 32'h00000000 /* 0x2764 */;
            2522: data_o = 32'h00000000 /* 0x2768 */;
            2523: data_o = 32'h00000000 /* 0x276c */;
            2524: data_o = 32'h00000000 /* 0x2770 */;
            2525: data_o = 32'h00000000 /* 0x2774 */;
            2526: data_o = 32'h00000000 /* 0x2778 */;
            2527: data_o = 32'h00000000 /* 0x277c */;
            2528: data_o = 32'h00000000 /* 0x2780 */;
            2529: data_o = 32'h00000000 /* 0x2784 */;
            2530: data_o = 32'h00000000 /* 0x2788 */;
            2531: data_o = 32'h00000000 /* 0x278c */;
            2532: data_o = 32'h00000000 /* 0x2790 */;
            2533: data_o = 32'h00000000 /* 0x2794 */;
            2534: data_o = 32'h00000000 /* 0x2798 */;
            2535: data_o = 32'h00000000 /* 0x279c */;
            2536: data_o = 32'h00000000 /* 0x27a0 */;
            2537: data_o = 32'h00000000 /* 0x27a4 */;
            2538: data_o = 32'h00000000 /* 0x27a8 */;
            2539: data_o = 32'h00000000 /* 0x27ac */;
            2540: data_o = 32'h00000000 /* 0x27b0 */;
            2541: data_o = 32'h00000000 /* 0x27b4 */;
            2542: data_o = 32'h00000000 /* 0x27b8 */;
            2543: data_o = 32'h00000000 /* 0x27bc */;
            2544: data_o = 32'h00000000 /* 0x27c0 */;
            2545: data_o = 32'h00000000 /* 0x27c4 */;
            2546: data_o = 32'h00000000 /* 0x27c8 */;
            2547: data_o = 32'h00000000 /* 0x27cc */;
            2548: data_o = 32'h00000000 /* 0x27d0 */;
            2549: data_o = 32'h00000000 /* 0x27d4 */;
            2550: data_o = 32'h00000000 /* 0x27d8 */;
            2551: data_o = 32'h00000000 /* 0x27dc */;
            2552: data_o = 32'h00000000 /* 0x27e0 */;
            2553: data_o = 32'h00000000 /* 0x27e4 */;
            2554: data_o = 32'h00000000 /* 0x27e8 */;
            2555: data_o = 32'h00000000 /* 0x27ec */;
            2556: data_o = 32'h00000000 /* 0x27f0 */;
            2557: data_o = 32'h00000000 /* 0x27f4 */;
            2558: data_o = 32'h00000000 /* 0x27f8 */;
            2559: data_o = 32'h00000000 /* 0x27fc */;
            2560: data_o = 32'h00000000 /* 0x2800 */;
            2561: data_o = 32'h00000000 /* 0x2804 */;
            2562: data_o = 32'h00000000 /* 0x2808 */;
            2563: data_o = 32'h00000000 /* 0x280c */;
            2564: data_o = 32'h00000000 /* 0x2810 */;
            2565: data_o = 32'h00000000 /* 0x2814 */;
            2566: data_o = 32'h00000000 /* 0x2818 */;
            2567: data_o = 32'h00000000 /* 0x281c */;
            2568: data_o = 32'h00000000 /* 0x2820 */;
            2569: data_o = 32'h00000000 /* 0x2824 */;
            2570: data_o = 32'h00000000 /* 0x2828 */;
            2571: data_o = 32'h00000000 /* 0x282c */;
            2572: data_o = 32'h00000000 /* 0x2830 */;
            2573: data_o = 32'h00000000 /* 0x2834 */;
            2574: data_o = 32'h00000000 /* 0x2838 */;
            2575: data_o = 32'h00000000 /* 0x283c */;
            2576: data_o = 32'h00000000 /* 0x2840 */;
            2577: data_o = 32'h00000000 /* 0x2844 */;
            2578: data_o = 32'h00000000 /* 0x2848 */;
            2579: data_o = 32'h00000000 /* 0x284c */;
            2580: data_o = 32'h00000000 /* 0x2850 */;
            2581: data_o = 32'h00000000 /* 0x2854 */;
            2582: data_o = 32'h00000000 /* 0x2858 */;
            2583: data_o = 32'h00000000 /* 0x285c */;
            2584: data_o = 32'h00000000 /* 0x2860 */;
            2585: data_o = 32'h00000000 /* 0x2864 */;
            2586: data_o = 32'h00000000 /* 0x2868 */;
            2587: data_o = 32'h00000000 /* 0x286c */;
            2588: data_o = 32'h00000000 /* 0x2870 */;
            2589: data_o = 32'h00000000 /* 0x2874 */;
            2590: data_o = 32'h00000000 /* 0x2878 */;
            2591: data_o = 32'h00000000 /* 0x287c */;
            2592: data_o = 32'h00000000 /* 0x2880 */;
            2593: data_o = 32'h00000000 /* 0x2884 */;
            2594: data_o = 32'h00000000 /* 0x2888 */;
            2595: data_o = 32'h00000000 /* 0x288c */;
            2596: data_o = 32'h00000000 /* 0x2890 */;
            2597: data_o = 32'h00000000 /* 0x2894 */;
            2598: data_o = 32'h00000000 /* 0x2898 */;
            2599: data_o = 32'h00000000 /* 0x289c */;
            2600: data_o = 32'h00000000 /* 0x28a0 */;
            2601: data_o = 32'h00000000 /* 0x28a4 */;
            2602: data_o = 32'h00000000 /* 0x28a8 */;
            2603: data_o = 32'h00000000 /* 0x28ac */;
            2604: data_o = 32'h00000000 /* 0x28b0 */;
            2605: data_o = 32'h00000000 /* 0x28b4 */;
            2606: data_o = 32'h00000000 /* 0x28b8 */;
            2607: data_o = 32'h00000000 /* 0x28bc */;
            2608: data_o = 32'h00000000 /* 0x28c0 */;
            2609: data_o = 32'h00000000 /* 0x28c4 */;
            2610: data_o = 32'h00000000 /* 0x28c8 */;
            2611: data_o = 32'h00000000 /* 0x28cc */;
            2612: data_o = 32'h00000000 /* 0x28d0 */;
            2613: data_o = 32'h00000000 /* 0x28d4 */;
            2614: data_o = 32'h00000000 /* 0x28d8 */;
            2615: data_o = 32'h00000000 /* 0x28dc */;
            2616: data_o = 32'h00000000 /* 0x28e0 */;
            2617: data_o = 32'h00000000 /* 0x28e4 */;
            2618: data_o = 32'h00000000 /* 0x28e8 */;
            2619: data_o = 32'h00000000 /* 0x28ec */;
            2620: data_o = 32'h00000000 /* 0x28f0 */;
            2621: data_o = 32'h00000000 /* 0x28f4 */;
            2622: data_o = 32'h00000000 /* 0x28f8 */;
            2623: data_o = 32'h00000000 /* 0x28fc */;
            2624: data_o = 32'h00000000 /* 0x2900 */;
            2625: data_o = 32'h00000000 /* 0x2904 */;
            2626: data_o = 32'h00000000 /* 0x2908 */;
            2627: data_o = 32'h00000000 /* 0x290c */;
            2628: data_o = 32'h00000000 /* 0x2910 */;
            2629: data_o = 32'h00000000 /* 0x2914 */;
            2630: data_o = 32'h00000000 /* 0x2918 */;
            2631: data_o = 32'h00000000 /* 0x291c */;
            2632: data_o = 32'h00000000 /* 0x2920 */;
            2633: data_o = 32'h00000000 /* 0x2924 */;
            2634: data_o = 32'h00000000 /* 0x2928 */;
            2635: data_o = 32'h00000000 /* 0x292c */;
            2636: data_o = 32'h00000000 /* 0x2930 */;
            2637: data_o = 32'h00000000 /* 0x2934 */;
            2638: data_o = 32'h00000000 /* 0x2938 */;
            2639: data_o = 32'h00000000 /* 0x293c */;
            2640: data_o = 32'h00000000 /* 0x2940 */;
            2641: data_o = 32'h00000000 /* 0x2944 */;
            2642: data_o = 32'h00000000 /* 0x2948 */;
            2643: data_o = 32'h00000000 /* 0x294c */;
            2644: data_o = 32'h00000000 /* 0x2950 */;
            2645: data_o = 32'h00000000 /* 0x2954 */;
            2646: data_o = 32'h00000000 /* 0x2958 */;
            2647: data_o = 32'h00000000 /* 0x295c */;
            2648: data_o = 32'h00000000 /* 0x2960 */;
            2649: data_o = 32'h00000000 /* 0x2964 */;
            2650: data_o = 32'h00000000 /* 0x2968 */;
            2651: data_o = 32'h00000000 /* 0x296c */;
            2652: data_o = 32'h00000000 /* 0x2970 */;
            2653: data_o = 32'h00000000 /* 0x2974 */;
            2654: data_o = 32'h00000000 /* 0x2978 */;
            2655: data_o = 32'h00000000 /* 0x297c */;
            2656: data_o = 32'h00000000 /* 0x2980 */;
            2657: data_o = 32'h00000000 /* 0x2984 */;
            2658: data_o = 32'h00000000 /* 0x2988 */;
            2659: data_o = 32'h00000000 /* 0x298c */;
            2660: data_o = 32'h00000000 /* 0x2990 */;
            2661: data_o = 32'h00000000 /* 0x2994 */;
            2662: data_o = 32'h00000000 /* 0x2998 */;
            2663: data_o = 32'h00000000 /* 0x299c */;
            2664: data_o = 32'h00000000 /* 0x29a0 */;
            2665: data_o = 32'h00000000 /* 0x29a4 */;
            2666: data_o = 32'h00000000 /* 0x29a8 */;
            2667: data_o = 32'h00000000 /* 0x29ac */;
            2668: data_o = 32'h00000000 /* 0x29b0 */;
            2669: data_o = 32'h00000000 /* 0x29b4 */;
            2670: data_o = 32'h00000000 /* 0x29b8 */;
            2671: data_o = 32'h00000000 /* 0x29bc */;
            2672: data_o = 32'h00000000 /* 0x29c0 */;
            2673: data_o = 32'h00000000 /* 0x29c4 */;
            2674: data_o = 32'h00000000 /* 0x29c8 */;
            2675: data_o = 32'h00000000 /* 0x29cc */;
            2676: data_o = 32'h00000000 /* 0x29d0 */;
            2677: data_o = 32'h00000000 /* 0x29d4 */;
            2678: data_o = 32'h00000000 /* 0x29d8 */;
            2679: data_o = 32'h00000000 /* 0x29dc */;
            2680: data_o = 32'h00000000 /* 0x29e0 */;
            2681: data_o = 32'h00000000 /* 0x29e4 */;
            2682: data_o = 32'h00000000 /* 0x29e8 */;
            2683: data_o = 32'h00000000 /* 0x29ec */;
            2684: data_o = 32'h00000000 /* 0x29f0 */;
            2685: data_o = 32'h00000000 /* 0x29f4 */;
            2686: data_o = 32'h00000000 /* 0x29f8 */;
            2687: data_o = 32'h00000000 /* 0x29fc */;
            2688: data_o = 32'h00000000 /* 0x2a00 */;
            2689: data_o = 32'h00000000 /* 0x2a04 */;
            2690: data_o = 32'h00000000 /* 0x2a08 */;
            2691: data_o = 32'h00000000 /* 0x2a0c */;
            2692: data_o = 32'h00000000 /* 0x2a10 */;
            2693: data_o = 32'h00000000 /* 0x2a14 */;
            2694: data_o = 32'h00000000 /* 0x2a18 */;
            2695: data_o = 32'h00000000 /* 0x2a1c */;
            2696: data_o = 32'h00000000 /* 0x2a20 */;
            2697: data_o = 32'h00000000 /* 0x2a24 */;
            2698: data_o = 32'h00000000 /* 0x2a28 */;
            2699: data_o = 32'h00000000 /* 0x2a2c */;
            2700: data_o = 32'h00000000 /* 0x2a30 */;
            2701: data_o = 32'h00000000 /* 0x2a34 */;
            2702: data_o = 32'h00000000 /* 0x2a38 */;
            2703: data_o = 32'h00000000 /* 0x2a3c */;
            2704: data_o = 32'h00000000 /* 0x2a40 */;
            2705: data_o = 32'h00000000 /* 0x2a44 */;
            2706: data_o = 32'h00000000 /* 0x2a48 */;
            2707: data_o = 32'h00000000 /* 0x2a4c */;
            2708: data_o = 32'h00000000 /* 0x2a50 */;
            2709: data_o = 32'h00000000 /* 0x2a54 */;
            2710: data_o = 32'h00000000 /* 0x2a58 */;
            2711: data_o = 32'h00000000 /* 0x2a5c */;
            2712: data_o = 32'h00000000 /* 0x2a60 */;
            2713: data_o = 32'h00000000 /* 0x2a64 */;
            2714: data_o = 32'h00000000 /* 0x2a68 */;
            2715: data_o = 32'h00000000 /* 0x2a6c */;
            2716: data_o = 32'h00000000 /* 0x2a70 */;
            2717: data_o = 32'h00000000 /* 0x2a74 */;
            2718: data_o = 32'h00000000 /* 0x2a78 */;
            2719: data_o = 32'h00000000 /* 0x2a7c */;
            2720: data_o = 32'h00000000 /* 0x2a80 */;
            2721: data_o = 32'h00000000 /* 0x2a84 */;
            2722: data_o = 32'h00000000 /* 0x2a88 */;
            2723: data_o = 32'h00000000 /* 0x2a8c */;
            2724: data_o = 32'h00000000 /* 0x2a90 */;
            2725: data_o = 32'h00000000 /* 0x2a94 */;
            2726: data_o = 32'h00000000 /* 0x2a98 */;
            2727: data_o = 32'h00000000 /* 0x2a9c */;
            2728: data_o = 32'h00000000 /* 0x2aa0 */;
            2729: data_o = 32'h00000000 /* 0x2aa4 */;
            2730: data_o = 32'h00000000 /* 0x2aa8 */;
            2731: data_o = 32'h00000000 /* 0x2aac */;
            2732: data_o = 32'h00000000 /* 0x2ab0 */;
            2733: data_o = 32'h00000000 /* 0x2ab4 */;
            2734: data_o = 32'h00000000 /* 0x2ab8 */;
            2735: data_o = 32'h00000000 /* 0x2abc */;
            2736: data_o = 32'h00000000 /* 0x2ac0 */;
            2737: data_o = 32'h00000000 /* 0x2ac4 */;
            2738: data_o = 32'h00000000 /* 0x2ac8 */;
            2739: data_o = 32'h00000000 /* 0x2acc */;
            2740: data_o = 32'h00000000 /* 0x2ad0 */;
            2741: data_o = 32'h00000000 /* 0x2ad4 */;
            2742: data_o = 32'h00000000 /* 0x2ad8 */;
            2743: data_o = 32'h00000000 /* 0x2adc */;
            2744: data_o = 32'h00000000 /* 0x2ae0 */;
            2745: data_o = 32'h00000000 /* 0x2ae4 */;
            2746: data_o = 32'h00000000 /* 0x2ae8 */;
            2747: data_o = 32'h00000000 /* 0x2aec */;
            2748: data_o = 32'h00000000 /* 0x2af0 */;
            2749: data_o = 32'h00000000 /* 0x2af4 */;
            2750: data_o = 32'h00000000 /* 0x2af8 */;
            2751: data_o = 32'h00000000 /* 0x2afc */;
            2752: data_o = 32'h00000000 /* 0x2b00 */;
            2753: data_o = 32'h00000000 /* 0x2b04 */;
            2754: data_o = 32'h00000000 /* 0x2b08 */;
            2755: data_o = 32'h00000000 /* 0x2b0c */;
            2756: data_o = 32'h00000000 /* 0x2b10 */;
            2757: data_o = 32'h00000000 /* 0x2b14 */;
            2758: data_o = 32'h00000000 /* 0x2b18 */;
            2759: data_o = 32'h00000000 /* 0x2b1c */;
            2760: data_o = 32'h00000000 /* 0x2b20 */;
            2761: data_o = 32'h00000000 /* 0x2b24 */;
            2762: data_o = 32'h00000000 /* 0x2b28 */;
            2763: data_o = 32'h00000000 /* 0x2b2c */;
            2764: data_o = 32'h00000000 /* 0x2b30 */;
            2765: data_o = 32'h00000000 /* 0x2b34 */;
            2766: data_o = 32'h00000000 /* 0x2b38 */;
            2767: data_o = 32'h00000000 /* 0x2b3c */;
            2768: data_o = 32'h00000000 /* 0x2b40 */;
            2769: data_o = 32'h00000000 /* 0x2b44 */;
            2770: data_o = 32'h00000000 /* 0x2b48 */;
            2771: data_o = 32'h00000000 /* 0x2b4c */;
            2772: data_o = 32'h00000000 /* 0x2b50 */;
            2773: data_o = 32'h00000000 /* 0x2b54 */;
            2774: data_o = 32'h00000000 /* 0x2b58 */;
            2775: data_o = 32'h00000000 /* 0x2b5c */;
            2776: data_o = 32'h00000000 /* 0x2b60 */;
            2777: data_o = 32'h00000000 /* 0x2b64 */;
            2778: data_o = 32'h00000000 /* 0x2b68 */;
            2779: data_o = 32'h00000000 /* 0x2b6c */;
            2780: data_o = 32'h00000000 /* 0x2b70 */;
            2781: data_o = 32'h00000000 /* 0x2b74 */;
            2782: data_o = 32'h00000000 /* 0x2b78 */;
            2783: data_o = 32'h00000000 /* 0x2b7c */;
            2784: data_o = 32'h00000000 /* 0x2b80 */;
            2785: data_o = 32'h00000000 /* 0x2b84 */;
            2786: data_o = 32'h00000000 /* 0x2b88 */;
            2787: data_o = 32'h00000000 /* 0x2b8c */;
            2788: data_o = 32'h00000000 /* 0x2b90 */;
            2789: data_o = 32'h00000000 /* 0x2b94 */;
            2790: data_o = 32'h00000000 /* 0x2b98 */;
            2791: data_o = 32'h00000000 /* 0x2b9c */;
            2792: data_o = 32'h00000000 /* 0x2ba0 */;
            2793: data_o = 32'h00000000 /* 0x2ba4 */;
            2794: data_o = 32'h00000000 /* 0x2ba8 */;
            2795: data_o = 32'h00000000 /* 0x2bac */;
            2796: data_o = 32'h00000000 /* 0x2bb0 */;
            2797: data_o = 32'h00000000 /* 0x2bb4 */;
            2798: data_o = 32'h00000000 /* 0x2bb8 */;
            2799: data_o = 32'h00000000 /* 0x2bbc */;
            2800: data_o = 32'h00000000 /* 0x2bc0 */;
            2801: data_o = 32'h00000000 /* 0x2bc4 */;
            2802: data_o = 32'h00000000 /* 0x2bc8 */;
            2803: data_o = 32'h00000000 /* 0x2bcc */;
            2804: data_o = 32'h00000000 /* 0x2bd0 */;
            2805: data_o = 32'h00000000 /* 0x2bd4 */;
            2806: data_o = 32'h00000000 /* 0x2bd8 */;
            2807: data_o = 32'h00000000 /* 0x2bdc */;
            2808: data_o = 32'h00000000 /* 0x2be0 */;
            2809: data_o = 32'h00000000 /* 0x2be4 */;
            2810: data_o = 32'h00000000 /* 0x2be8 */;
            2811: data_o = 32'h00000000 /* 0x2bec */;
            2812: data_o = 32'h00000000 /* 0x2bf0 */;
            2813: data_o = 32'h00000000 /* 0x2bf4 */;
            2814: data_o = 32'h00000000 /* 0x2bf8 */;
            2815: data_o = 32'h00000000 /* 0x2bfc */;
            2816: data_o = 32'h00000000 /* 0x2c00 */;
            2817: data_o = 32'h00000000 /* 0x2c04 */;
            2818: data_o = 32'h00000000 /* 0x2c08 */;
            2819: data_o = 32'h00000000 /* 0x2c0c */;
            2820: data_o = 32'h00000000 /* 0x2c10 */;
            2821: data_o = 32'h00000000 /* 0x2c14 */;
            2822: data_o = 32'h00000000 /* 0x2c18 */;
            2823: data_o = 32'h00000000 /* 0x2c1c */;
            2824: data_o = 32'h00000000 /* 0x2c20 */;
            2825: data_o = 32'h00000000 /* 0x2c24 */;
            2826: data_o = 32'h00000000 /* 0x2c28 */;
            2827: data_o = 32'h00000000 /* 0x2c2c */;
            2828: data_o = 32'h00000000 /* 0x2c30 */;
            2829: data_o = 32'h00000000 /* 0x2c34 */;
            2830: data_o = 32'h00000000 /* 0x2c38 */;
            2831: data_o = 32'h00000000 /* 0x2c3c */;
            2832: data_o = 32'h00000000 /* 0x2c40 */;
            2833: data_o = 32'h00000000 /* 0x2c44 */;
            2834: data_o = 32'h00000000 /* 0x2c48 */;
            2835: data_o = 32'h00000000 /* 0x2c4c */;
            2836: data_o = 32'h00000000 /* 0x2c50 */;
            2837: data_o = 32'h00000000 /* 0x2c54 */;
            2838: data_o = 32'h00000000 /* 0x2c58 */;
            2839: data_o = 32'h00000000 /* 0x2c5c */;
            2840: data_o = 32'h00000000 /* 0x2c60 */;
            2841: data_o = 32'h00000000 /* 0x2c64 */;
            2842: data_o = 32'h00000000 /* 0x2c68 */;
            2843: data_o = 32'h00000000 /* 0x2c6c */;
            2844: data_o = 32'h00000000 /* 0x2c70 */;
            2845: data_o = 32'h00000000 /* 0x2c74 */;
            2846: data_o = 32'h00000000 /* 0x2c78 */;
            2847: data_o = 32'h00000000 /* 0x2c7c */;
            2848: data_o = 32'h00000000 /* 0x2c80 */;
            2849: data_o = 32'h00000000 /* 0x2c84 */;
            2850: data_o = 32'h00000000 /* 0x2c88 */;
            2851: data_o = 32'h00000000 /* 0x2c8c */;
            2852: data_o = 32'h00000000 /* 0x2c90 */;
            2853: data_o = 32'h00000000 /* 0x2c94 */;
            2854: data_o = 32'h00000000 /* 0x2c98 */;
            2855: data_o = 32'h00000000 /* 0x2c9c */;
            2856: data_o = 32'h00000000 /* 0x2ca0 */;
            2857: data_o = 32'h00000000 /* 0x2ca4 */;
            2858: data_o = 32'h00000000 /* 0x2ca8 */;
            2859: data_o = 32'h00000000 /* 0x2cac */;
            2860: data_o = 32'h00000000 /* 0x2cb0 */;
            2861: data_o = 32'h00000000 /* 0x2cb4 */;
            2862: data_o = 32'h00000000 /* 0x2cb8 */;
            2863: data_o = 32'h00000000 /* 0x2cbc */;
            2864: data_o = 32'h00000000 /* 0x2cc0 */;
            2865: data_o = 32'h00000000 /* 0x2cc4 */;
            2866: data_o = 32'h00000000 /* 0x2cc8 */;
            2867: data_o = 32'h00000000 /* 0x2ccc */;
            2868: data_o = 32'h00000000 /* 0x2cd0 */;
            2869: data_o = 32'h00000000 /* 0x2cd4 */;
            2870: data_o = 32'h00000000 /* 0x2cd8 */;
            2871: data_o = 32'h00000000 /* 0x2cdc */;
            2872: data_o = 32'h00000000 /* 0x2ce0 */;
            2873: data_o = 32'h00000000 /* 0x2ce4 */;
            2874: data_o = 32'h00000000 /* 0x2ce8 */;
            2875: data_o = 32'h00000000 /* 0x2cec */;
            2876: data_o = 32'h00000000 /* 0x2cf0 */;
            2877: data_o = 32'h00000000 /* 0x2cf4 */;
            2878: data_o = 32'h00000000 /* 0x2cf8 */;
            2879: data_o = 32'h00000000 /* 0x2cfc */;
            2880: data_o = 32'h00000000 /* 0x2d00 */;
            2881: data_o = 32'h00000000 /* 0x2d04 */;
            2882: data_o = 32'h00000000 /* 0x2d08 */;
            2883: data_o = 32'h00000000 /* 0x2d0c */;
            2884: data_o = 32'h00000000 /* 0x2d10 */;
            2885: data_o = 32'h00000000 /* 0x2d14 */;
            2886: data_o = 32'h00000000 /* 0x2d18 */;
            2887: data_o = 32'h00000000 /* 0x2d1c */;
            2888: data_o = 32'h00000000 /* 0x2d20 */;
            2889: data_o = 32'h00000000 /* 0x2d24 */;
            2890: data_o = 32'h00000000 /* 0x2d28 */;
            2891: data_o = 32'h00000000 /* 0x2d2c */;
            2892: data_o = 32'h00000000 /* 0x2d30 */;
            2893: data_o = 32'h00000000 /* 0x2d34 */;
            2894: data_o = 32'h00000000 /* 0x2d38 */;
            2895: data_o = 32'h00000000 /* 0x2d3c */;
            2896: data_o = 32'h00000000 /* 0x2d40 */;
            2897: data_o = 32'h00000000 /* 0x2d44 */;
            2898: data_o = 32'h00000000 /* 0x2d48 */;
            2899: data_o = 32'h00000000 /* 0x2d4c */;
            2900: data_o = 32'h00000000 /* 0x2d50 */;
            2901: data_o = 32'h00000000 /* 0x2d54 */;
            2902: data_o = 32'h00000000 /* 0x2d58 */;
            2903: data_o = 32'h00000000 /* 0x2d5c */;
            2904: data_o = 32'h00000000 /* 0x2d60 */;
            2905: data_o = 32'h00000000 /* 0x2d64 */;
            2906: data_o = 32'h00000000 /* 0x2d68 */;
            2907: data_o = 32'h00000000 /* 0x2d6c */;
            2908: data_o = 32'h00000000 /* 0x2d70 */;
            2909: data_o = 32'h00000000 /* 0x2d74 */;
            2910: data_o = 32'h00000000 /* 0x2d78 */;
            2911: data_o = 32'h00000000 /* 0x2d7c */;
            2912: data_o = 32'h00000000 /* 0x2d80 */;
            2913: data_o = 32'h00000000 /* 0x2d84 */;
            2914: data_o = 32'h00000000 /* 0x2d88 */;
            2915: data_o = 32'h00000000 /* 0x2d8c */;
            2916: data_o = 32'h00000000 /* 0x2d90 */;
            2917: data_o = 32'h00000000 /* 0x2d94 */;
            2918: data_o = 32'h00000000 /* 0x2d98 */;
            2919: data_o = 32'h00000000 /* 0x2d9c */;
            2920: data_o = 32'h00000000 /* 0x2da0 */;
            2921: data_o = 32'h00000000 /* 0x2da4 */;
            2922: data_o = 32'h00000000 /* 0x2da8 */;
            2923: data_o = 32'h00000000 /* 0x2dac */;
            2924: data_o = 32'h00000000 /* 0x2db0 */;
            2925: data_o = 32'h00000000 /* 0x2db4 */;
            2926: data_o = 32'h00000000 /* 0x2db8 */;
            2927: data_o = 32'h00000000 /* 0x2dbc */;
            2928: data_o = 32'h00000000 /* 0x2dc0 */;
            2929: data_o = 32'h00000000 /* 0x2dc4 */;
            2930: data_o = 32'h00000000 /* 0x2dc8 */;
            2931: data_o = 32'h00000000 /* 0x2dcc */;
            2932: data_o = 32'h00000000 /* 0x2dd0 */;
            2933: data_o = 32'h00000000 /* 0x2dd4 */;
            2934: data_o = 32'h00000000 /* 0x2dd8 */;
            2935: data_o = 32'h00000000 /* 0x2ddc */;
            2936: data_o = 32'h00000000 /* 0x2de0 */;
            2937: data_o = 32'h00000000 /* 0x2de4 */;
            2938: data_o = 32'h00000000 /* 0x2de8 */;
            2939: data_o = 32'h00000000 /* 0x2dec */;
            2940: data_o = 32'h00000000 /* 0x2df0 */;
            2941: data_o = 32'h00000000 /* 0x2df4 */;
            2942: data_o = 32'h00000000 /* 0x2df8 */;
            2943: data_o = 32'h00000000 /* 0x2dfc */;
            2944: data_o = 32'h00000000 /* 0x2e00 */;
            2945: data_o = 32'h00000000 /* 0x2e04 */;
            2946: data_o = 32'h00000000 /* 0x2e08 */;
            2947: data_o = 32'h00000000 /* 0x2e0c */;
            2948: data_o = 32'h00000000 /* 0x2e10 */;
            2949: data_o = 32'h00000000 /* 0x2e14 */;
            2950: data_o = 32'h00000000 /* 0x2e18 */;
            2951: data_o = 32'h00000000 /* 0x2e1c */;
            2952: data_o = 32'h00000000 /* 0x2e20 */;
            2953: data_o = 32'h00000000 /* 0x2e24 */;
            2954: data_o = 32'h00000000 /* 0x2e28 */;
            2955: data_o = 32'h00000000 /* 0x2e2c */;
            2956: data_o = 32'h00000000 /* 0x2e30 */;
            2957: data_o = 32'h00000000 /* 0x2e34 */;
            2958: data_o = 32'h00000000 /* 0x2e38 */;
            2959: data_o = 32'h00000000 /* 0x2e3c */;
            2960: data_o = 32'h00000000 /* 0x2e40 */;
            2961: data_o = 32'h00000000 /* 0x2e44 */;
            2962: data_o = 32'h00000000 /* 0x2e48 */;
            2963: data_o = 32'h00000000 /* 0x2e4c */;
            2964: data_o = 32'h00000000 /* 0x2e50 */;
            2965: data_o = 32'h00000000 /* 0x2e54 */;
            2966: data_o = 32'h00000000 /* 0x2e58 */;
            2967: data_o = 32'h00000000 /* 0x2e5c */;
            2968: data_o = 32'h00000000 /* 0x2e60 */;
            2969: data_o = 32'h00000000 /* 0x2e64 */;
            2970: data_o = 32'h00000000 /* 0x2e68 */;
            2971: data_o = 32'h00000000 /* 0x2e6c */;
            2972: data_o = 32'h00000000 /* 0x2e70 */;
            2973: data_o = 32'h00000000 /* 0x2e74 */;
            2974: data_o = 32'h00000000 /* 0x2e78 */;
            2975: data_o = 32'h00000000 /* 0x2e7c */;
            2976: data_o = 32'h00000000 /* 0x2e80 */;
            2977: data_o = 32'h00000000 /* 0x2e84 */;
            2978: data_o = 32'h00000000 /* 0x2e88 */;
            2979: data_o = 32'h00000000 /* 0x2e8c */;
            2980: data_o = 32'h00000000 /* 0x2e90 */;
            2981: data_o = 32'h00000000 /* 0x2e94 */;
            2982: data_o = 32'h00000000 /* 0x2e98 */;
            2983: data_o = 32'h00000000 /* 0x2e9c */;
            2984: data_o = 32'h00000000 /* 0x2ea0 */;
            2985: data_o = 32'h00000000 /* 0x2ea4 */;
            2986: data_o = 32'h00000000 /* 0x2ea8 */;
            2987: data_o = 32'h00000000 /* 0x2eac */;
            2988: data_o = 32'h00000000 /* 0x2eb0 */;
            2989: data_o = 32'h00000000 /* 0x2eb4 */;
            2990: data_o = 32'h00000000 /* 0x2eb8 */;
            2991: data_o = 32'h00000000 /* 0x2ebc */;
            2992: data_o = 32'h00000000 /* 0x2ec0 */;
            2993: data_o = 32'h00000000 /* 0x2ec4 */;
            2994: data_o = 32'h00000000 /* 0x2ec8 */;
            2995: data_o = 32'h00000000 /* 0x2ecc */;
            2996: data_o = 32'h00000000 /* 0x2ed0 */;
            2997: data_o = 32'h00000000 /* 0x2ed4 */;
            2998: data_o = 32'h00000000 /* 0x2ed8 */;
            2999: data_o = 32'h00000000 /* 0x2edc */;
            3000: data_o = 32'h00000000 /* 0x2ee0 */;
            3001: data_o = 32'h00000000 /* 0x2ee4 */;
            3002: data_o = 32'h00000000 /* 0x2ee8 */;
            3003: data_o = 32'h00000000 /* 0x2eec */;
            3004: data_o = 32'h00000000 /* 0x2ef0 */;
            3005: data_o = 32'h00000000 /* 0x2ef4 */;
            3006: data_o = 32'h00000000 /* 0x2ef8 */;
            3007: data_o = 32'h00000000 /* 0x2efc */;
            3008: data_o = 32'h00000000 /* 0x2f00 */;
            3009: data_o = 32'h00000000 /* 0x2f04 */;
            3010: data_o = 32'h00000000 /* 0x2f08 */;
            3011: data_o = 32'h00000000 /* 0x2f0c */;
            3012: data_o = 32'h00000000 /* 0x2f10 */;
            3013: data_o = 32'h00000000 /* 0x2f14 */;
            3014: data_o = 32'h00000000 /* 0x2f18 */;
            3015: data_o = 32'h00000000 /* 0x2f1c */;
            3016: data_o = 32'h00000000 /* 0x2f20 */;
            3017: data_o = 32'h00000000 /* 0x2f24 */;
            3018: data_o = 32'h00000000 /* 0x2f28 */;
            3019: data_o = 32'h00000000 /* 0x2f2c */;
            3020: data_o = 32'h00000000 /* 0x2f30 */;
            3021: data_o = 32'h00000000 /* 0x2f34 */;
            3022: data_o = 32'h00000000 /* 0x2f38 */;
            3023: data_o = 32'h00000000 /* 0x2f3c */;
            3024: data_o = 32'h00000000 /* 0x2f40 */;
            3025: data_o = 32'h00000000 /* 0x2f44 */;
            3026: data_o = 32'h00000000 /* 0x2f48 */;
            3027: data_o = 32'h00000000 /* 0x2f4c */;
            3028: data_o = 32'h00000000 /* 0x2f50 */;
            3029: data_o = 32'h00000000 /* 0x2f54 */;
            3030: data_o = 32'h00000000 /* 0x2f58 */;
            3031: data_o = 32'h00000000 /* 0x2f5c */;
            3032: data_o = 32'h00000000 /* 0x2f60 */;
            3033: data_o = 32'h00000000 /* 0x2f64 */;
            3034: data_o = 32'h00000000 /* 0x2f68 */;
            3035: data_o = 32'h00000000 /* 0x2f6c */;
            3036: data_o = 32'h00000000 /* 0x2f70 */;
            3037: data_o = 32'h00000000 /* 0x2f74 */;
            3038: data_o = 32'h00000000 /* 0x2f78 */;
            3039: data_o = 32'h00000000 /* 0x2f7c */;
            3040: data_o = 32'h00000000 /* 0x2f80 */;
            3041: data_o = 32'h00000000 /* 0x2f84 */;
            3042: data_o = 32'h00000000 /* 0x2f88 */;
            3043: data_o = 32'h00000000 /* 0x2f8c */;
            3044: data_o = 32'h00000000 /* 0x2f90 */;
            3045: data_o = 32'h00000000 /* 0x2f94 */;
            3046: data_o = 32'h00000000 /* 0x2f98 */;
            3047: data_o = 32'h00000000 /* 0x2f9c */;
            3048: data_o = 32'h00000000 /* 0x2fa0 */;
            3049: data_o = 32'h00000000 /* 0x2fa4 */;
            3050: data_o = 32'h00000000 /* 0x2fa8 */;
            3051: data_o = 32'h00000000 /* 0x2fac */;
            3052: data_o = 32'h00000000 /* 0x2fb0 */;
            3053: data_o = 32'h00000000 /* 0x2fb4 */;
            3054: data_o = 32'h00000000 /* 0x2fb8 */;
            3055: data_o = 32'h00000000 /* 0x2fbc */;
            3056: data_o = 32'h00000000 /* 0x2fc0 */;
            3057: data_o = 32'h00000000 /* 0x2fc4 */;
            3058: data_o = 32'h00000000 /* 0x2fc8 */;
            3059: data_o = 32'h00000000 /* 0x2fcc */;
            3060: data_o = 32'h00000000 /* 0x2fd0 */;
            3061: data_o = 32'h00000000 /* 0x2fd4 */;
            3062: data_o = 32'h00000000 /* 0x2fd8 */;
            3063: data_o = 32'h00000000 /* 0x2fdc */;
            3064: data_o = 32'h00000000 /* 0x2fe0 */;
            3065: data_o = 32'h00000000 /* 0x2fe4 */;
            3066: data_o = 32'h00000000 /* 0x2fe8 */;
            3067: data_o = 32'h00000000 /* 0x2fec */;
            3068: data_o = 32'h00000000 /* 0x2ff0 */;
            3069: data_o = 32'h00000000 /* 0x2ff4 */;
            3070: data_o = 32'h00000000 /* 0x2ff8 */;
            3071: data_o = 32'h00000000 /* 0x2ffc */;
            3072: data_o = 32'h00000000 /* 0x3000 */;
            3073: data_o = 32'h00000000 /* 0x3004 */;
            3074: data_o = 32'h00000000 /* 0x3008 */;
            3075: data_o = 32'h00000000 /* 0x300c */;
            3076: data_o = 32'h00000000 /* 0x3010 */;
            3077: data_o = 32'h00000000 /* 0x3014 */;
            3078: data_o = 32'h00000000 /* 0x3018 */;
            3079: data_o = 32'h00000000 /* 0x301c */;
            3080: data_o = 32'h00000000 /* 0x3020 */;
            3081: data_o = 32'h00000000 /* 0x3024 */;
            3082: data_o = 32'h00000000 /* 0x3028 */;
            3083: data_o = 32'h00000000 /* 0x302c */;
            3084: data_o = 32'h00000000 /* 0x3030 */;
            3085: data_o = 32'h00000000 /* 0x3034 */;
            3086: data_o = 32'h00000000 /* 0x3038 */;
            3087: data_o = 32'h00000000 /* 0x303c */;
            3088: data_o = 32'h00000000 /* 0x3040 */;
            3089: data_o = 32'h00000000 /* 0x3044 */;
            3090: data_o = 32'h00000000 /* 0x3048 */;
            3091: data_o = 32'h00000000 /* 0x304c */;
            3092: data_o = 32'h00000000 /* 0x3050 */;
            3093: data_o = 32'h00000000 /* 0x3054 */;
            3094: data_o = 32'h00000000 /* 0x3058 */;
            3095: data_o = 32'h00000000 /* 0x305c */;
            3096: data_o = 32'h00000000 /* 0x3060 */;
            3097: data_o = 32'h00000000 /* 0x3064 */;
            3098: data_o = 32'h00000000 /* 0x3068 */;
            3099: data_o = 32'h00000000 /* 0x306c */;
            3100: data_o = 32'h00000000 /* 0x3070 */;
            3101: data_o = 32'h00000000 /* 0x3074 */;
            3102: data_o = 32'h00000000 /* 0x3078 */;
            3103: data_o = 32'h00000000 /* 0x307c */;
            3104: data_o = 32'h00000000 /* 0x3080 */;
            3105: data_o = 32'h00000000 /* 0x3084 */;
            3106: data_o = 32'h00000000 /* 0x3088 */;
            3107: data_o = 32'h00000000 /* 0x308c */;
            3108: data_o = 32'h00000000 /* 0x3090 */;
            3109: data_o = 32'h00000000 /* 0x3094 */;
            3110: data_o = 32'h00000000 /* 0x3098 */;
            3111: data_o = 32'h00000000 /* 0x309c */;
            3112: data_o = 32'h00000000 /* 0x30a0 */;
            3113: data_o = 32'h00000000 /* 0x30a4 */;
            3114: data_o = 32'h00000000 /* 0x30a8 */;
            3115: data_o = 32'h00000000 /* 0x30ac */;
            3116: data_o = 32'h00000000 /* 0x30b0 */;
            3117: data_o = 32'h00000000 /* 0x30b4 */;
            3118: data_o = 32'h00000000 /* 0x30b8 */;
            3119: data_o = 32'h00000000 /* 0x30bc */;
            3120: data_o = 32'h00000000 /* 0x30c0 */;
            3121: data_o = 32'h00000000 /* 0x30c4 */;
            3122: data_o = 32'h00000000 /* 0x30c8 */;
            3123: data_o = 32'h00000000 /* 0x30cc */;
            3124: data_o = 32'h00000000 /* 0x30d0 */;
            3125: data_o = 32'h00000000 /* 0x30d4 */;
            3126: data_o = 32'h00000000 /* 0x30d8 */;
            3127: data_o = 32'h00000000 /* 0x30dc */;
            3128: data_o = 32'h00000000 /* 0x30e0 */;
            3129: data_o = 32'h00000000 /* 0x30e4 */;
            3130: data_o = 32'h00000000 /* 0x30e8 */;
            3131: data_o = 32'h00000000 /* 0x30ec */;
            3132: data_o = 32'h00000000 /* 0x30f0 */;
            3133: data_o = 32'h00000000 /* 0x30f4 */;
            3134: data_o = 32'h00000000 /* 0x30f8 */;
            3135: data_o = 32'h00000000 /* 0x30fc */;
            3136: data_o = 32'h00000000 /* 0x3100 */;
            3137: data_o = 32'h00000000 /* 0x3104 */;
            3138: data_o = 32'h00000000 /* 0x3108 */;
            3139: data_o = 32'h00000000 /* 0x310c */;
            3140: data_o = 32'h00000000 /* 0x3110 */;
            3141: data_o = 32'h00000000 /* 0x3114 */;
            3142: data_o = 32'h00000000 /* 0x3118 */;
            3143: data_o = 32'h00000000 /* 0x311c */;
            3144: data_o = 32'h00000000 /* 0x3120 */;
            3145: data_o = 32'h00000000 /* 0x3124 */;
            3146: data_o = 32'h00000000 /* 0x3128 */;
            3147: data_o = 32'h00000000 /* 0x312c */;
            3148: data_o = 32'h00000000 /* 0x3130 */;
            3149: data_o = 32'h00000000 /* 0x3134 */;
            3150: data_o = 32'h00000000 /* 0x3138 */;
            3151: data_o = 32'h00000000 /* 0x313c */;
            3152: data_o = 32'h00000000 /* 0x3140 */;
            3153: data_o = 32'h00000000 /* 0x3144 */;
            3154: data_o = 32'h00000000 /* 0x3148 */;
            3155: data_o = 32'h00000000 /* 0x314c */;
            3156: data_o = 32'h00000000 /* 0x3150 */;
            3157: data_o = 32'h00000000 /* 0x3154 */;
            3158: data_o = 32'h00000000 /* 0x3158 */;
            3159: data_o = 32'h00000000 /* 0x315c */;
            3160: data_o = 32'h00000000 /* 0x3160 */;
            3161: data_o = 32'h00000000 /* 0x3164 */;
            3162: data_o = 32'h00000000 /* 0x3168 */;
            3163: data_o = 32'h00000000 /* 0x316c */;
            3164: data_o = 32'h00000000 /* 0x3170 */;
            3165: data_o = 32'h00000000 /* 0x3174 */;
            3166: data_o = 32'h00000000 /* 0x3178 */;
            3167: data_o = 32'h00000000 /* 0x317c */;
            3168: data_o = 32'h00000000 /* 0x3180 */;
            3169: data_o = 32'h00000000 /* 0x3184 */;
            3170: data_o = 32'h00000000 /* 0x3188 */;
            3171: data_o = 32'h00000000 /* 0x318c */;
            3172: data_o = 32'h00000000 /* 0x3190 */;
            3173: data_o = 32'h00000000 /* 0x3194 */;
            3174: data_o = 32'h00000000 /* 0x3198 */;
            3175: data_o = 32'h00000000 /* 0x319c */;
            3176: data_o = 32'h00000000 /* 0x31a0 */;
            3177: data_o = 32'h00000000 /* 0x31a4 */;
            3178: data_o = 32'h00000000 /* 0x31a8 */;
            3179: data_o = 32'h00000000 /* 0x31ac */;
            3180: data_o = 32'h00000000 /* 0x31b0 */;
            3181: data_o = 32'h00000000 /* 0x31b4 */;
            3182: data_o = 32'h00000000 /* 0x31b8 */;
            3183: data_o = 32'h00000000 /* 0x31bc */;
            3184: data_o = 32'h00000000 /* 0x31c0 */;
            3185: data_o = 32'h00000000 /* 0x31c4 */;
            3186: data_o = 32'h00000000 /* 0x31c8 */;
            3187: data_o = 32'h00000000 /* 0x31cc */;
            3188: data_o = 32'h00000000 /* 0x31d0 */;
            3189: data_o = 32'h00000000 /* 0x31d4 */;
            3190: data_o = 32'h00000000 /* 0x31d8 */;
            3191: data_o = 32'h00000000 /* 0x31dc */;
            3192: data_o = 32'h00000000 /* 0x31e0 */;
            3193: data_o = 32'h00000000 /* 0x31e4 */;
            3194: data_o = 32'h00000000 /* 0x31e8 */;
            3195: data_o = 32'h00000000 /* 0x31ec */;
            3196: data_o = 32'h00000000 /* 0x31f0 */;
            3197: data_o = 32'h00000000 /* 0x31f4 */;
            3198: data_o = 32'h00000000 /* 0x31f8 */;
            3199: data_o = 32'h00000000 /* 0x31fc */;
            3200: data_o = 32'h00000000 /* 0x3200 */;
            3201: data_o = 32'h00000000 /* 0x3204 */;
            3202: data_o = 32'h00000000 /* 0x3208 */;
            3203: data_o = 32'h00000000 /* 0x320c */;
            3204: data_o = 32'h00000000 /* 0x3210 */;
            3205: data_o = 32'h00000000 /* 0x3214 */;
            3206: data_o = 32'h00000000 /* 0x3218 */;
            3207: data_o = 32'h00000000 /* 0x321c */;
            3208: data_o = 32'h00000000 /* 0x3220 */;
            3209: data_o = 32'h00000000 /* 0x3224 */;
            3210: data_o = 32'h00000000 /* 0x3228 */;
            3211: data_o = 32'h00000000 /* 0x322c */;
            3212: data_o = 32'h00000000 /* 0x3230 */;
            3213: data_o = 32'h00000000 /* 0x3234 */;
            3214: data_o = 32'h00000000 /* 0x3238 */;
            3215: data_o = 32'h00000000 /* 0x323c */;
            3216: data_o = 32'h00000000 /* 0x3240 */;
            3217: data_o = 32'h00000000 /* 0x3244 */;
            3218: data_o = 32'h00000000 /* 0x3248 */;
            3219: data_o = 32'h00000000 /* 0x324c */;
            3220: data_o = 32'h00000000 /* 0x3250 */;
            3221: data_o = 32'h00000000 /* 0x3254 */;
            3222: data_o = 32'h00000000 /* 0x3258 */;
            3223: data_o = 32'h00000000 /* 0x325c */;
            3224: data_o = 32'h00000000 /* 0x3260 */;
            3225: data_o = 32'h00000000 /* 0x3264 */;
            3226: data_o = 32'h00000000 /* 0x3268 */;
            3227: data_o = 32'h00000000 /* 0x326c */;
            3228: data_o = 32'h00000000 /* 0x3270 */;
            3229: data_o = 32'h00000000 /* 0x3274 */;
            3230: data_o = 32'h00000000 /* 0x3278 */;
            3231: data_o = 32'h00000000 /* 0x327c */;
            3232: data_o = 32'h00000000 /* 0x3280 */;
            3233: data_o = 32'h00000000 /* 0x3284 */;
            3234: data_o = 32'h00000000 /* 0x3288 */;
            3235: data_o = 32'h00000000 /* 0x328c */;
            3236: data_o = 32'h00000000 /* 0x3290 */;
            3237: data_o = 32'h00000000 /* 0x3294 */;
            3238: data_o = 32'h00000000 /* 0x3298 */;
            3239: data_o = 32'h00000000 /* 0x329c */;
            3240: data_o = 32'h00000000 /* 0x32a0 */;
            3241: data_o = 32'h00000000 /* 0x32a4 */;
            3242: data_o = 32'h00000000 /* 0x32a8 */;
            3243: data_o = 32'h00000000 /* 0x32ac */;
            3244: data_o = 32'h00000000 /* 0x32b0 */;
            3245: data_o = 32'h00000000 /* 0x32b4 */;
            3246: data_o = 32'h00000000 /* 0x32b8 */;
            3247: data_o = 32'h00000000 /* 0x32bc */;
            3248: data_o = 32'h00000000 /* 0x32c0 */;
            3249: data_o = 32'h00000000 /* 0x32c4 */;
            3250: data_o = 32'h00000000 /* 0x32c8 */;
            3251: data_o = 32'h00000000 /* 0x32cc */;
            3252: data_o = 32'h00000000 /* 0x32d0 */;
            3253: data_o = 32'h00000000 /* 0x32d4 */;
            3254: data_o = 32'h00000000 /* 0x32d8 */;
            3255: data_o = 32'h00000000 /* 0x32dc */;
            3256: data_o = 32'h00000000 /* 0x32e0 */;
            3257: data_o = 32'h00000000 /* 0x32e4 */;
            3258: data_o = 32'h00000000 /* 0x32e8 */;
            3259: data_o = 32'h00000000 /* 0x32ec */;
            3260: data_o = 32'h00000000 /* 0x32f0 */;
            3261: data_o = 32'h00000000 /* 0x32f4 */;
            3262: data_o = 32'h00000000 /* 0x32f8 */;
            3263: data_o = 32'h00000000 /* 0x32fc */;
            3264: data_o = 32'h00000000 /* 0x3300 */;
            3265: data_o = 32'h00000000 /* 0x3304 */;
            3266: data_o = 32'h00000000 /* 0x3308 */;
            3267: data_o = 32'h00000000 /* 0x330c */;
            3268: data_o = 32'h00000000 /* 0x3310 */;
            3269: data_o = 32'h00000000 /* 0x3314 */;
            3270: data_o = 32'h00000000 /* 0x3318 */;
            3271: data_o = 32'h00000000 /* 0x331c */;
            3272: data_o = 32'h00000000 /* 0x3320 */;
            3273: data_o = 32'h00000000 /* 0x3324 */;
            3274: data_o = 32'h00000000 /* 0x3328 */;
            3275: data_o = 32'h00000000 /* 0x332c */;
            3276: data_o = 32'h00000000 /* 0x3330 */;
            3277: data_o = 32'h00000000 /* 0x3334 */;
            3278: data_o = 32'h00000000 /* 0x3338 */;
            3279: data_o = 32'h00000000 /* 0x333c */;
            3280: data_o = 32'h00000000 /* 0x3340 */;
            3281: data_o = 32'h00000000 /* 0x3344 */;
            3282: data_o = 32'h00000000 /* 0x3348 */;
            3283: data_o = 32'h00000000 /* 0x334c */;
            3284: data_o = 32'h00000000 /* 0x3350 */;
            3285: data_o = 32'h00000000 /* 0x3354 */;
            3286: data_o = 32'h00000000 /* 0x3358 */;
            3287: data_o = 32'h00000000 /* 0x335c */;
            3288: data_o = 32'h00000000 /* 0x3360 */;
            3289: data_o = 32'h00000000 /* 0x3364 */;
            3290: data_o = 32'h00000000 /* 0x3368 */;
            3291: data_o = 32'h00000000 /* 0x336c */;
            3292: data_o = 32'h00000000 /* 0x3370 */;
            3293: data_o = 32'h00000000 /* 0x3374 */;
            3294: data_o = 32'h00000000 /* 0x3378 */;
            3295: data_o = 32'h00000000 /* 0x337c */;
            3296: data_o = 32'h00000000 /* 0x3380 */;
            3297: data_o = 32'h00000000 /* 0x3384 */;
            3298: data_o = 32'h00000000 /* 0x3388 */;
            3299: data_o = 32'h00000000 /* 0x338c */;
            3300: data_o = 32'h00000000 /* 0x3390 */;
            3301: data_o = 32'h00000000 /* 0x3394 */;
            3302: data_o = 32'h00000000 /* 0x3398 */;
            3303: data_o = 32'h00000000 /* 0x339c */;
            3304: data_o = 32'h00000000 /* 0x33a0 */;
            3305: data_o = 32'h00000000 /* 0x33a4 */;
            3306: data_o = 32'h00000000 /* 0x33a8 */;
            3307: data_o = 32'h00000000 /* 0x33ac */;
            3308: data_o = 32'h00000000 /* 0x33b0 */;
            3309: data_o = 32'h00000000 /* 0x33b4 */;
            3310: data_o = 32'h00000000 /* 0x33b8 */;
            3311: data_o = 32'h00000000 /* 0x33bc */;
            3312: data_o = 32'h00000000 /* 0x33c0 */;
            3313: data_o = 32'h00000000 /* 0x33c4 */;
            3314: data_o = 32'h00000000 /* 0x33c8 */;
            3315: data_o = 32'h00000000 /* 0x33cc */;
            3316: data_o = 32'h00000000 /* 0x33d0 */;
            3317: data_o = 32'h00000000 /* 0x33d4 */;
            3318: data_o = 32'h00000000 /* 0x33d8 */;
            3319: data_o = 32'h00000000 /* 0x33dc */;
            3320: data_o = 32'h00000000 /* 0x33e0 */;
            3321: data_o = 32'h00000000 /* 0x33e4 */;
            3322: data_o = 32'h00000000 /* 0x33e8 */;
            3323: data_o = 32'h00000000 /* 0x33ec */;
            3324: data_o = 32'h00000000 /* 0x33f0 */;
            3325: data_o = 32'h00000000 /* 0x33f4 */;
            3326: data_o = 32'h00000000 /* 0x33f8 */;
            3327: data_o = 32'h00000000 /* 0x33fc */;
            3328: data_o = 32'h00000000 /* 0x3400 */;
            3329: data_o = 32'h00000000 /* 0x3404 */;
            3330: data_o = 32'h00000000 /* 0x3408 */;
            3331: data_o = 32'h00000000 /* 0x340c */;
            3332: data_o = 32'h00000000 /* 0x3410 */;
            3333: data_o = 32'h00000000 /* 0x3414 */;
            3334: data_o = 32'h00000000 /* 0x3418 */;
            3335: data_o = 32'h00000000 /* 0x341c */;
            3336: data_o = 32'h00000000 /* 0x3420 */;
            3337: data_o = 32'h00000000 /* 0x3424 */;
            3338: data_o = 32'h00000000 /* 0x3428 */;
            3339: data_o = 32'h00000000 /* 0x342c */;
            3340: data_o = 32'h00000000 /* 0x3430 */;
            3341: data_o = 32'h00000000 /* 0x3434 */;
            3342: data_o = 32'h00000000 /* 0x3438 */;
            3343: data_o = 32'h00000000 /* 0x343c */;
            3344: data_o = 32'h00000000 /* 0x3440 */;
            3345: data_o = 32'h00000000 /* 0x3444 */;
            3346: data_o = 32'h00000000 /* 0x3448 */;
            3347: data_o = 32'h00000000 /* 0x344c */;
            3348: data_o = 32'h00000000 /* 0x3450 */;
            3349: data_o = 32'h00000000 /* 0x3454 */;
            3350: data_o = 32'h00000000 /* 0x3458 */;
            3351: data_o = 32'h00000000 /* 0x345c */;
            3352: data_o = 32'h00000000 /* 0x3460 */;
            3353: data_o = 32'h00000000 /* 0x3464 */;
            3354: data_o = 32'h00000000 /* 0x3468 */;
            3355: data_o = 32'h00000000 /* 0x346c */;
            3356: data_o = 32'h00000000 /* 0x3470 */;
            3357: data_o = 32'h00000000 /* 0x3474 */;
            3358: data_o = 32'h00000000 /* 0x3478 */;
            3359: data_o = 32'h00000000 /* 0x347c */;
            3360: data_o = 32'h00000000 /* 0x3480 */;
            3361: data_o = 32'h00000000 /* 0x3484 */;
            3362: data_o = 32'h00000000 /* 0x3488 */;
            3363: data_o = 32'h00000000 /* 0x348c */;
            3364: data_o = 32'h00000000 /* 0x3490 */;
            3365: data_o = 32'h00000000 /* 0x3494 */;
            3366: data_o = 32'h00000000 /* 0x3498 */;
            3367: data_o = 32'h00000000 /* 0x349c */;
            3368: data_o = 32'h00000000 /* 0x34a0 */;
            3369: data_o = 32'h00000000 /* 0x34a4 */;
            3370: data_o = 32'h00000000 /* 0x34a8 */;
            3371: data_o = 32'h00000000 /* 0x34ac */;
            3372: data_o = 32'h00000000 /* 0x34b0 */;
            3373: data_o = 32'h00000000 /* 0x34b4 */;
            3374: data_o = 32'h00000000 /* 0x34b8 */;
            3375: data_o = 32'h00000000 /* 0x34bc */;
            3376: data_o = 32'h00000000 /* 0x34c0 */;
            3377: data_o = 32'h00000000 /* 0x34c4 */;
            3378: data_o = 32'h00000000 /* 0x34c8 */;
            3379: data_o = 32'h00000000 /* 0x34cc */;
            3380: data_o = 32'h00000000 /* 0x34d0 */;
            3381: data_o = 32'h00000000 /* 0x34d4 */;
            3382: data_o = 32'h00000000 /* 0x34d8 */;
            3383: data_o = 32'h00000000 /* 0x34dc */;
            3384: data_o = 32'h00000000 /* 0x34e0 */;
            3385: data_o = 32'h00000000 /* 0x34e4 */;
            3386: data_o = 32'h00000000 /* 0x34e8 */;
            3387: data_o = 32'h00000000 /* 0x34ec */;
            3388: data_o = 32'h00000000 /* 0x34f0 */;
            3389: data_o = 32'h00000000 /* 0x34f4 */;
            3390: data_o = 32'h00000000 /* 0x34f8 */;
            3391: data_o = 32'h00000000 /* 0x34fc */;
            3392: data_o = 32'h00000000 /* 0x3500 */;
            3393: data_o = 32'h00000000 /* 0x3504 */;
            3394: data_o = 32'h00000000 /* 0x3508 */;
            3395: data_o = 32'h00000000 /* 0x350c */;
            3396: data_o = 32'h00000000 /* 0x3510 */;
            3397: data_o = 32'h00000000 /* 0x3514 */;
            3398: data_o = 32'h00000000 /* 0x3518 */;
            3399: data_o = 32'h00000000 /* 0x351c */;
            3400: data_o = 32'h00000000 /* 0x3520 */;
            3401: data_o = 32'h00000000 /* 0x3524 */;
            3402: data_o = 32'h00000000 /* 0x3528 */;
            3403: data_o = 32'h00000000 /* 0x352c */;
            3404: data_o = 32'h00000000 /* 0x3530 */;
            3405: data_o = 32'h00000000 /* 0x3534 */;
            3406: data_o = 32'h00000000 /* 0x3538 */;
            3407: data_o = 32'h00000000 /* 0x353c */;
            3408: data_o = 32'h00000000 /* 0x3540 */;
            3409: data_o = 32'h00000000 /* 0x3544 */;
            3410: data_o = 32'h00000000 /* 0x3548 */;
            3411: data_o = 32'h00000000 /* 0x354c */;
            3412: data_o = 32'h00000000 /* 0x3550 */;
            3413: data_o = 32'h00000000 /* 0x3554 */;
            3414: data_o = 32'h00000000 /* 0x3558 */;
            3415: data_o = 32'h00000000 /* 0x355c */;
            3416: data_o = 32'h00000000 /* 0x3560 */;
            3417: data_o = 32'h00000000 /* 0x3564 */;
            3418: data_o = 32'h00000000 /* 0x3568 */;
            3419: data_o = 32'h00000000 /* 0x356c */;
            3420: data_o = 32'h00000000 /* 0x3570 */;
            3421: data_o = 32'h00000000 /* 0x3574 */;
            3422: data_o = 32'h00000000 /* 0x3578 */;
            3423: data_o = 32'h00000000 /* 0x357c */;
            3424: data_o = 32'h00000000 /* 0x3580 */;
            3425: data_o = 32'h00000000 /* 0x3584 */;
            3426: data_o = 32'h00000000 /* 0x3588 */;
            3427: data_o = 32'h00000000 /* 0x358c */;
            3428: data_o = 32'h00000000 /* 0x3590 */;
            3429: data_o = 32'h00000000 /* 0x3594 */;
            3430: data_o = 32'h00000000 /* 0x3598 */;
            3431: data_o = 32'h00000000 /* 0x359c */;
            3432: data_o = 32'h00000000 /* 0x35a0 */;
            3433: data_o = 32'h00000000 /* 0x35a4 */;
            3434: data_o = 32'h00000000 /* 0x35a8 */;
            3435: data_o = 32'h00000000 /* 0x35ac */;
            3436: data_o = 32'h00000000 /* 0x35b0 */;
            3437: data_o = 32'h00000000 /* 0x35b4 */;
            3438: data_o = 32'h00000000 /* 0x35b8 */;
            3439: data_o = 32'h00000000 /* 0x35bc */;
            3440: data_o = 32'h00000000 /* 0x35c0 */;
            3441: data_o = 32'h00000000 /* 0x35c4 */;
            3442: data_o = 32'h00000000 /* 0x35c8 */;
            3443: data_o = 32'h00000000 /* 0x35cc */;
            3444: data_o = 32'h00000000 /* 0x35d0 */;
            3445: data_o = 32'h00000000 /* 0x35d4 */;
            3446: data_o = 32'h00000000 /* 0x35d8 */;
            3447: data_o = 32'h00000000 /* 0x35dc */;
            3448: data_o = 32'h00000000 /* 0x35e0 */;
            3449: data_o = 32'h00000000 /* 0x35e4 */;
            3450: data_o = 32'h00000000 /* 0x35e8 */;
            3451: data_o = 32'h00000000 /* 0x35ec */;
            3452: data_o = 32'h00000000 /* 0x35f0 */;
            3453: data_o = 32'h00000000 /* 0x35f4 */;
            3454: data_o = 32'h00000000 /* 0x35f8 */;
            3455: data_o = 32'h00000000 /* 0x35fc */;
            3456: data_o = 32'h00000000 /* 0x3600 */;
            3457: data_o = 32'h00000000 /* 0x3604 */;
            3458: data_o = 32'h00000000 /* 0x3608 */;
            3459: data_o = 32'h00000000 /* 0x360c */;
            3460: data_o = 32'h00000000 /* 0x3610 */;
            3461: data_o = 32'h00000000 /* 0x3614 */;
            3462: data_o = 32'h00000000 /* 0x3618 */;
            3463: data_o = 32'h00000000 /* 0x361c */;
            3464: data_o = 32'h00000000 /* 0x3620 */;
            3465: data_o = 32'h00000000 /* 0x3624 */;
            3466: data_o = 32'h00000000 /* 0x3628 */;
            3467: data_o = 32'h00000000 /* 0x362c */;
            3468: data_o = 32'h00000000 /* 0x3630 */;
            3469: data_o = 32'h00000000 /* 0x3634 */;
            3470: data_o = 32'h00000000 /* 0x3638 */;
            3471: data_o = 32'h00000000 /* 0x363c */;
            3472: data_o = 32'h00000000 /* 0x3640 */;
            3473: data_o = 32'h00000000 /* 0x3644 */;
            3474: data_o = 32'h00000000 /* 0x3648 */;
            3475: data_o = 32'h00000000 /* 0x364c */;
            3476: data_o = 32'h00000000 /* 0x3650 */;
            3477: data_o = 32'h00000000 /* 0x3654 */;
            3478: data_o = 32'h00000000 /* 0x3658 */;
            3479: data_o = 32'h00000000 /* 0x365c */;
            3480: data_o = 32'h00000000 /* 0x3660 */;
            3481: data_o = 32'h00000000 /* 0x3664 */;
            3482: data_o = 32'h00000000 /* 0x3668 */;
            3483: data_o = 32'h00000000 /* 0x366c */;
            3484: data_o = 32'h00000000 /* 0x3670 */;
            3485: data_o = 32'h00000000 /* 0x3674 */;
            3486: data_o = 32'h00000000 /* 0x3678 */;
            3487: data_o = 32'h00000000 /* 0x367c */;
            3488: data_o = 32'h00000000 /* 0x3680 */;
            3489: data_o = 32'h00000000 /* 0x3684 */;
            3490: data_o = 32'h00000000 /* 0x3688 */;
            3491: data_o = 32'h00000000 /* 0x368c */;
            3492: data_o = 32'h00000000 /* 0x3690 */;
            3493: data_o = 32'h00000000 /* 0x3694 */;
            3494: data_o = 32'h00000000 /* 0x3698 */;
            3495: data_o = 32'h00000000 /* 0x369c */;
            3496: data_o = 32'h00000000 /* 0x36a0 */;
            3497: data_o = 32'h00000000 /* 0x36a4 */;
            3498: data_o = 32'h00000000 /* 0x36a8 */;
            3499: data_o = 32'h00000000 /* 0x36ac */;
            3500: data_o = 32'h00000000 /* 0x36b0 */;
            3501: data_o = 32'h00000000 /* 0x36b4 */;
            3502: data_o = 32'h00000000 /* 0x36b8 */;
            3503: data_o = 32'h00000000 /* 0x36bc */;
            3504: data_o = 32'h00000000 /* 0x36c0 */;
            3505: data_o = 32'h00000000 /* 0x36c4 */;
            3506: data_o = 32'h00000000 /* 0x36c8 */;
            3507: data_o = 32'h00000000 /* 0x36cc */;
            3508: data_o = 32'h00000000 /* 0x36d0 */;
            3509: data_o = 32'h00000000 /* 0x36d4 */;
            3510: data_o = 32'h00000000 /* 0x36d8 */;
            3511: data_o = 32'h00000000 /* 0x36dc */;
            3512: data_o = 32'h00000000 /* 0x36e0 */;
            3513: data_o = 32'h00000000 /* 0x36e4 */;
            3514: data_o = 32'h00000000 /* 0x36e8 */;
            3515: data_o = 32'h00000000 /* 0x36ec */;
            3516: data_o = 32'h00000000 /* 0x36f0 */;
            3517: data_o = 32'h00000000 /* 0x36f4 */;
            3518: data_o = 32'h00000000 /* 0x36f8 */;
            3519: data_o = 32'h00000000 /* 0x36fc */;
            3520: data_o = 32'h00000000 /* 0x3700 */;
            3521: data_o = 32'h00000000 /* 0x3704 */;
            3522: data_o = 32'h00000000 /* 0x3708 */;
            3523: data_o = 32'h00000000 /* 0x370c */;
            3524: data_o = 32'h00000000 /* 0x3710 */;
            3525: data_o = 32'h00000000 /* 0x3714 */;
            3526: data_o = 32'h00000000 /* 0x3718 */;
            3527: data_o = 32'h00000000 /* 0x371c */;
            3528: data_o = 32'h00000000 /* 0x3720 */;
            3529: data_o = 32'h00000000 /* 0x3724 */;
            3530: data_o = 32'h00000000 /* 0x3728 */;
            3531: data_o = 32'h00000000 /* 0x372c */;
            3532: data_o = 32'h00000000 /* 0x3730 */;
            3533: data_o = 32'h00000000 /* 0x3734 */;
            3534: data_o = 32'h00000000 /* 0x3738 */;
            3535: data_o = 32'h00000000 /* 0x373c */;
            3536: data_o = 32'h00000000 /* 0x3740 */;
            3537: data_o = 32'h00000000 /* 0x3744 */;
            3538: data_o = 32'h00000000 /* 0x3748 */;
            3539: data_o = 32'h00000000 /* 0x374c */;
            3540: data_o = 32'h00000000 /* 0x3750 */;
            3541: data_o = 32'h00000000 /* 0x3754 */;
            3542: data_o = 32'h00000000 /* 0x3758 */;
            3543: data_o = 32'h00000000 /* 0x375c */;
            3544: data_o = 32'h00000000 /* 0x3760 */;
            3545: data_o = 32'h00000000 /* 0x3764 */;
            3546: data_o = 32'h00000000 /* 0x3768 */;
            3547: data_o = 32'h00000000 /* 0x376c */;
            3548: data_o = 32'h00000000 /* 0x3770 */;
            3549: data_o = 32'h00000000 /* 0x3774 */;
            3550: data_o = 32'h00000000 /* 0x3778 */;
            3551: data_o = 32'h00000000 /* 0x377c */;
            3552: data_o = 32'h00000000 /* 0x3780 */;
            3553: data_o = 32'h00000000 /* 0x3784 */;
            3554: data_o = 32'h00000000 /* 0x3788 */;
            3555: data_o = 32'h00000000 /* 0x378c */;
            3556: data_o = 32'h00000000 /* 0x3790 */;
            3557: data_o = 32'h00000000 /* 0x3794 */;
            3558: data_o = 32'h00000000 /* 0x3798 */;
            3559: data_o = 32'h00000000 /* 0x379c */;
            3560: data_o = 32'h00000000 /* 0x37a0 */;
            3561: data_o = 32'h00000000 /* 0x37a4 */;
            3562: data_o = 32'h00000000 /* 0x37a8 */;
            3563: data_o = 32'h00000000 /* 0x37ac */;
            3564: data_o = 32'h00000000 /* 0x37b0 */;
            3565: data_o = 32'h00000000 /* 0x37b4 */;
            3566: data_o = 32'h00000000 /* 0x37b8 */;
            3567: data_o = 32'h00000000 /* 0x37bc */;
            3568: data_o = 32'h00000000 /* 0x37c0 */;
            3569: data_o = 32'h00000000 /* 0x37c4 */;
            3570: data_o = 32'h00000000 /* 0x37c8 */;
            3571: data_o = 32'h00000000 /* 0x37cc */;
            3572: data_o = 32'h00000000 /* 0x37d0 */;
            3573: data_o = 32'h00000000 /* 0x37d4 */;
            3574: data_o = 32'h00000000 /* 0x37d8 */;
            3575: data_o = 32'h00000000 /* 0x37dc */;
            3576: data_o = 32'h00000000 /* 0x37e0 */;
            3577: data_o = 32'h00000000 /* 0x37e4 */;
            3578: data_o = 32'h00000000 /* 0x37e8 */;
            3579: data_o = 32'h00000000 /* 0x37ec */;
            3580: data_o = 32'h00000000 /* 0x37f0 */;
            3581: data_o = 32'h00000000 /* 0x37f4 */;
            3582: data_o = 32'h00000000 /* 0x37f8 */;
            3583: data_o = 32'h00000000 /* 0x37fc */;
            3584: data_o = 32'h00000000 /* 0x3800 */;
            3585: data_o = 32'h00000000 /* 0x3804 */;
            3586: data_o = 32'h00000000 /* 0x3808 */;
            3587: data_o = 32'h00000000 /* 0x380c */;
            3588: data_o = 32'h00000000 /* 0x3810 */;
            3589: data_o = 32'h00000000 /* 0x3814 */;
            3590: data_o = 32'h00000000 /* 0x3818 */;
            3591: data_o = 32'h00000000 /* 0x381c */;
            3592: data_o = 32'h00000000 /* 0x3820 */;
            3593: data_o = 32'h00000000 /* 0x3824 */;
            3594: data_o = 32'h00000000 /* 0x3828 */;
            3595: data_o = 32'h00000000 /* 0x382c */;
            3596: data_o = 32'h00000000 /* 0x3830 */;
            3597: data_o = 32'h00000000 /* 0x3834 */;
            3598: data_o = 32'h00000000 /* 0x3838 */;
            3599: data_o = 32'h00000000 /* 0x383c */;
            3600: data_o = 32'h00000000 /* 0x3840 */;
            3601: data_o = 32'h00000000 /* 0x3844 */;
            3602: data_o = 32'h00000000 /* 0x3848 */;
            3603: data_o = 32'h00000000 /* 0x384c */;
            3604: data_o = 32'h00000000 /* 0x3850 */;
            3605: data_o = 32'h00000000 /* 0x3854 */;
            3606: data_o = 32'h00000000 /* 0x3858 */;
            3607: data_o = 32'h00000000 /* 0x385c */;
            3608: data_o = 32'h00000000 /* 0x3860 */;
            3609: data_o = 32'h00000000 /* 0x3864 */;
            3610: data_o = 32'h00000000 /* 0x3868 */;
            3611: data_o = 32'h00000000 /* 0x386c */;
            3612: data_o = 32'h00000000 /* 0x3870 */;
            3613: data_o = 32'h00000000 /* 0x3874 */;
            3614: data_o = 32'h00000000 /* 0x3878 */;
            3615: data_o = 32'h00000000 /* 0x387c */;
            3616: data_o = 32'h00000000 /* 0x3880 */;
            3617: data_o = 32'h00000000 /* 0x3884 */;
            3618: data_o = 32'h00000000 /* 0x3888 */;
            3619: data_o = 32'h00000000 /* 0x388c */;
            3620: data_o = 32'h00000000 /* 0x3890 */;
            3621: data_o = 32'h00000000 /* 0x3894 */;
            3622: data_o = 32'h00000000 /* 0x3898 */;
            3623: data_o = 32'h00000000 /* 0x389c */;
            3624: data_o = 32'h00000000 /* 0x38a0 */;
            3625: data_o = 32'h00000000 /* 0x38a4 */;
            3626: data_o = 32'h00000000 /* 0x38a8 */;
            3627: data_o = 32'h00000000 /* 0x38ac */;
            3628: data_o = 32'h00000000 /* 0x38b0 */;
            3629: data_o = 32'h00000000 /* 0x38b4 */;
            3630: data_o = 32'h00000000 /* 0x38b8 */;
            3631: data_o = 32'h00000000 /* 0x38bc */;
            3632: data_o = 32'h00000000 /* 0x38c0 */;
            3633: data_o = 32'h00000000 /* 0x38c4 */;
            3634: data_o = 32'h00000000 /* 0x38c8 */;
            3635: data_o = 32'h00000000 /* 0x38cc */;
            3636: data_o = 32'h00000000 /* 0x38d0 */;
            3637: data_o = 32'h00000000 /* 0x38d4 */;
            3638: data_o = 32'h00000000 /* 0x38d8 */;
            3639: data_o = 32'h00000000 /* 0x38dc */;
            3640: data_o = 32'h00000000 /* 0x38e0 */;
            3641: data_o = 32'h00000000 /* 0x38e4 */;
            3642: data_o = 32'h00000000 /* 0x38e8 */;
            3643: data_o = 32'h00000000 /* 0x38ec */;
            3644: data_o = 32'h00000000 /* 0x38f0 */;
            3645: data_o = 32'h00000000 /* 0x38f4 */;
            3646: data_o = 32'h00000000 /* 0x38f8 */;
            3647: data_o = 32'h00000000 /* 0x38fc */;
            3648: data_o = 32'h00000000 /* 0x3900 */;
            3649: data_o = 32'h00000000 /* 0x3904 */;
            3650: data_o = 32'h00000000 /* 0x3908 */;
            3651: data_o = 32'h00000000 /* 0x390c */;
            3652: data_o = 32'h00000000 /* 0x3910 */;
            3653: data_o = 32'h00000000 /* 0x3914 */;
            3654: data_o = 32'h00000000 /* 0x3918 */;
            3655: data_o = 32'h00000000 /* 0x391c */;
            3656: data_o = 32'h00000000 /* 0x3920 */;
            3657: data_o = 32'h00000000 /* 0x3924 */;
            3658: data_o = 32'h00000000 /* 0x3928 */;
            3659: data_o = 32'h00000000 /* 0x392c */;
            3660: data_o = 32'h00000000 /* 0x3930 */;
            3661: data_o = 32'h00000000 /* 0x3934 */;
            3662: data_o = 32'h00000000 /* 0x3938 */;
            3663: data_o = 32'h00000000 /* 0x393c */;
            3664: data_o = 32'h00000000 /* 0x3940 */;
            3665: data_o = 32'h00000000 /* 0x3944 */;
            3666: data_o = 32'h00000000 /* 0x3948 */;
            3667: data_o = 32'h00000000 /* 0x394c */;
            3668: data_o = 32'h00000000 /* 0x3950 */;
            3669: data_o = 32'h00000000 /* 0x3954 */;
            3670: data_o = 32'h00000000 /* 0x3958 */;
            3671: data_o = 32'h00000000 /* 0x395c */;
            3672: data_o = 32'h00000000 /* 0x3960 */;
            3673: data_o = 32'h00000000 /* 0x3964 */;
            3674: data_o = 32'h00000000 /* 0x3968 */;
            3675: data_o = 32'h00000000 /* 0x396c */;
            3676: data_o = 32'h00000000 /* 0x3970 */;
            3677: data_o = 32'h00000000 /* 0x3974 */;
            3678: data_o = 32'h00000000 /* 0x3978 */;
            3679: data_o = 32'h00000000 /* 0x397c */;
            3680: data_o = 32'h00000000 /* 0x3980 */;
            3681: data_o = 32'h00000000 /* 0x3984 */;
            3682: data_o = 32'h00000000 /* 0x3988 */;
            3683: data_o = 32'h00000000 /* 0x398c */;
            3684: data_o = 32'h00000000 /* 0x3990 */;
            3685: data_o = 32'h00000000 /* 0x3994 */;
            3686: data_o = 32'h00000000 /* 0x3998 */;
            3687: data_o = 32'h00000000 /* 0x399c */;
            3688: data_o = 32'h00000000 /* 0x39a0 */;
            3689: data_o = 32'h00000000 /* 0x39a4 */;
            3690: data_o = 32'h00000000 /* 0x39a8 */;
            3691: data_o = 32'h00000000 /* 0x39ac */;
            3692: data_o = 32'h00000000 /* 0x39b0 */;
            3693: data_o = 32'h00000000 /* 0x39b4 */;
            3694: data_o = 32'h00000000 /* 0x39b8 */;
            3695: data_o = 32'h00000000 /* 0x39bc */;
            3696: data_o = 32'h00000000 /* 0x39c0 */;
            3697: data_o = 32'h00000000 /* 0x39c4 */;
            3698: data_o = 32'h00000000 /* 0x39c8 */;
            3699: data_o = 32'h00000000 /* 0x39cc */;
            3700: data_o = 32'h00000000 /* 0x39d0 */;
            3701: data_o = 32'h00000000 /* 0x39d4 */;
            3702: data_o = 32'h00000000 /* 0x39d8 */;
            3703: data_o = 32'h00000000 /* 0x39dc */;
            3704: data_o = 32'h00000000 /* 0x39e0 */;
            3705: data_o = 32'h00000000 /* 0x39e4 */;
            3706: data_o = 32'h00000000 /* 0x39e8 */;
            3707: data_o = 32'h00000000 /* 0x39ec */;
            3708: data_o = 32'h00000000 /* 0x39f0 */;
            3709: data_o = 32'h00000000 /* 0x39f4 */;
            3710: data_o = 32'h00000000 /* 0x39f8 */;
            3711: data_o = 32'h00000000 /* 0x39fc */;
            3712: data_o = 32'h00000000 /* 0x3a00 */;
            3713: data_o = 32'h00000000 /* 0x3a04 */;
            3714: data_o = 32'h00000000 /* 0x3a08 */;
            3715: data_o = 32'h00000000 /* 0x3a0c */;
            3716: data_o = 32'h00000000 /* 0x3a10 */;
            3717: data_o = 32'h00000000 /* 0x3a14 */;
            3718: data_o = 32'h00000000 /* 0x3a18 */;
            3719: data_o = 32'h00000000 /* 0x3a1c */;
            3720: data_o = 32'h00000000 /* 0x3a20 */;
            3721: data_o = 32'h00000000 /* 0x3a24 */;
            3722: data_o = 32'h00000000 /* 0x3a28 */;
            3723: data_o = 32'h00000000 /* 0x3a2c */;
            3724: data_o = 32'h00000000 /* 0x3a30 */;
            3725: data_o = 32'h00000000 /* 0x3a34 */;
            3726: data_o = 32'h00000000 /* 0x3a38 */;
            3727: data_o = 32'h00000000 /* 0x3a3c */;
            3728: data_o = 32'h00000000 /* 0x3a40 */;
            3729: data_o = 32'h00000000 /* 0x3a44 */;
            3730: data_o = 32'h00000000 /* 0x3a48 */;
            3731: data_o = 32'h00000000 /* 0x3a4c */;
            3732: data_o = 32'h00000000 /* 0x3a50 */;
            3733: data_o = 32'h00000000 /* 0x3a54 */;
            3734: data_o = 32'h00000000 /* 0x3a58 */;
            3735: data_o = 32'h00000000 /* 0x3a5c */;
            3736: data_o = 32'h00000000 /* 0x3a60 */;
            3737: data_o = 32'h00000000 /* 0x3a64 */;
            3738: data_o = 32'h00000000 /* 0x3a68 */;
            3739: data_o = 32'h00000000 /* 0x3a6c */;
            3740: data_o = 32'h00000000 /* 0x3a70 */;
            3741: data_o = 32'h00000000 /* 0x3a74 */;
            3742: data_o = 32'h00000000 /* 0x3a78 */;
            3743: data_o = 32'h00000000 /* 0x3a7c */;
            3744: data_o = 32'h00000000 /* 0x3a80 */;
            3745: data_o = 32'h00000000 /* 0x3a84 */;
            3746: data_o = 32'h00000000 /* 0x3a88 */;
            3747: data_o = 32'h00000000 /* 0x3a8c */;
            3748: data_o = 32'h00000000 /* 0x3a90 */;
            3749: data_o = 32'h00000000 /* 0x3a94 */;
            3750: data_o = 32'h00000000 /* 0x3a98 */;
            3751: data_o = 32'h00000000 /* 0x3a9c */;
            3752: data_o = 32'h00000000 /* 0x3aa0 */;
            3753: data_o = 32'h00000000 /* 0x3aa4 */;
            3754: data_o = 32'h00000000 /* 0x3aa8 */;
            3755: data_o = 32'h00000000 /* 0x3aac */;
            3756: data_o = 32'h00000000 /* 0x3ab0 */;
            3757: data_o = 32'h00000000 /* 0x3ab4 */;
            3758: data_o = 32'h00000000 /* 0x3ab8 */;
            3759: data_o = 32'h00000000 /* 0x3abc */;
            3760: data_o = 32'h00000000 /* 0x3ac0 */;
            3761: data_o = 32'h00000000 /* 0x3ac4 */;
            3762: data_o = 32'h00000000 /* 0x3ac8 */;
            3763: data_o = 32'h00000000 /* 0x3acc */;
            3764: data_o = 32'h00000000 /* 0x3ad0 */;
            3765: data_o = 32'h00000000 /* 0x3ad4 */;
            3766: data_o = 32'h00000000 /* 0x3ad8 */;
            3767: data_o = 32'h00000000 /* 0x3adc */;
            3768: data_o = 32'h00000000 /* 0x3ae0 */;
            3769: data_o = 32'h00000000 /* 0x3ae4 */;
            3770: data_o = 32'h00000000 /* 0x3ae8 */;
            3771: data_o = 32'h00000000 /* 0x3aec */;
            3772: data_o = 32'h00000000 /* 0x3af0 */;
            3773: data_o = 32'h00000000 /* 0x3af4 */;
            3774: data_o = 32'h00000000 /* 0x3af8 */;
            3775: data_o = 32'h00000000 /* 0x3afc */;
            3776: data_o = 32'h00000000 /* 0x3b00 */;
            3777: data_o = 32'h00000000 /* 0x3b04 */;
            3778: data_o = 32'h00000000 /* 0x3b08 */;
            3779: data_o = 32'h00000000 /* 0x3b0c */;
            3780: data_o = 32'h00000000 /* 0x3b10 */;
            3781: data_o = 32'h00000000 /* 0x3b14 */;
            3782: data_o = 32'h00000000 /* 0x3b18 */;
            3783: data_o = 32'h00000000 /* 0x3b1c */;
            3784: data_o = 32'h00000000 /* 0x3b20 */;
            3785: data_o = 32'h00000000 /* 0x3b24 */;
            3786: data_o = 32'h00000000 /* 0x3b28 */;
            3787: data_o = 32'h00000000 /* 0x3b2c */;
            3788: data_o = 32'h00000000 /* 0x3b30 */;
            3789: data_o = 32'h00000000 /* 0x3b34 */;
            3790: data_o = 32'h00000000 /* 0x3b38 */;
            3791: data_o = 32'h00000000 /* 0x3b3c */;
            3792: data_o = 32'h00000000 /* 0x3b40 */;
            3793: data_o = 32'h00000000 /* 0x3b44 */;
            3794: data_o = 32'h00000000 /* 0x3b48 */;
            3795: data_o = 32'h00000000 /* 0x3b4c */;
            3796: data_o = 32'h00000000 /* 0x3b50 */;
            3797: data_o = 32'h00000000 /* 0x3b54 */;
            3798: data_o = 32'h00000000 /* 0x3b58 */;
            3799: data_o = 32'h00000000 /* 0x3b5c */;
            3800: data_o = 32'h00000000 /* 0x3b60 */;
            3801: data_o = 32'h00000000 /* 0x3b64 */;
            3802: data_o = 32'h00000000 /* 0x3b68 */;
            3803: data_o = 32'h00000000 /* 0x3b6c */;
            3804: data_o = 32'h00000000 /* 0x3b70 */;
            3805: data_o = 32'h00000000 /* 0x3b74 */;
            3806: data_o = 32'h00000000 /* 0x3b78 */;
            3807: data_o = 32'h00000000 /* 0x3b7c */;
            3808: data_o = 32'h00000000 /* 0x3b80 */;
            3809: data_o = 32'h00000000 /* 0x3b84 */;
            3810: data_o = 32'h00000000 /* 0x3b88 */;
            3811: data_o = 32'h00000000 /* 0x3b8c */;
            3812: data_o = 32'h00000000 /* 0x3b90 */;
            3813: data_o = 32'h00000000 /* 0x3b94 */;
            3814: data_o = 32'h00000000 /* 0x3b98 */;
            3815: data_o = 32'h00000000 /* 0x3b9c */;
            3816: data_o = 32'h00000000 /* 0x3ba0 */;
            3817: data_o = 32'h00000000 /* 0x3ba4 */;
            3818: data_o = 32'h00000000 /* 0x3ba8 */;
            3819: data_o = 32'h00000000 /* 0x3bac */;
            3820: data_o = 32'h00000000 /* 0x3bb0 */;
            3821: data_o = 32'h00000000 /* 0x3bb4 */;
            3822: data_o = 32'h00000000 /* 0x3bb8 */;
            3823: data_o = 32'h00000000 /* 0x3bbc */;
            3824: data_o = 32'h00000000 /* 0x3bc0 */;
            3825: data_o = 32'h00000000 /* 0x3bc4 */;
            3826: data_o = 32'h00000000 /* 0x3bc8 */;
            3827: data_o = 32'h00000000 /* 0x3bcc */;
            3828: data_o = 32'h00000000 /* 0x3bd0 */;
            3829: data_o = 32'h00000000 /* 0x3bd4 */;
            3830: data_o = 32'h00000000 /* 0x3bd8 */;
            3831: data_o = 32'h00000000 /* 0x3bdc */;
            3832: data_o = 32'h00000000 /* 0x3be0 */;
            3833: data_o = 32'h00000000 /* 0x3be4 */;
            3834: data_o = 32'h00000000 /* 0x3be8 */;
            3835: data_o = 32'h00000000 /* 0x3bec */;
            3836: data_o = 32'h00000000 /* 0x3bf0 */;
            3837: data_o = 32'h00000000 /* 0x3bf4 */;
            3838: data_o = 32'h00000000 /* 0x3bf8 */;
            3839: data_o = 32'h00000000 /* 0x3bfc */;
            3840: data_o = 32'h00000000 /* 0x3c00 */;
            3841: data_o = 32'h00000000 /* 0x3c04 */;
            3842: data_o = 32'h00000000 /* 0x3c08 */;
            3843: data_o = 32'h00000000 /* 0x3c0c */;
            3844: data_o = 32'h00000000 /* 0x3c10 */;
            3845: data_o = 32'h00000000 /* 0x3c14 */;
            3846: data_o = 32'h00000000 /* 0x3c18 */;
            3847: data_o = 32'h00000000 /* 0x3c1c */;
            3848: data_o = 32'h00000000 /* 0x3c20 */;
            3849: data_o = 32'h00000000 /* 0x3c24 */;
            3850: data_o = 32'h00000000 /* 0x3c28 */;
            3851: data_o = 32'h00000000 /* 0x3c2c */;
            3852: data_o = 32'h00000000 /* 0x3c30 */;
            3853: data_o = 32'h00000000 /* 0x3c34 */;
            3854: data_o = 32'h00000000 /* 0x3c38 */;
            3855: data_o = 32'h00000000 /* 0x3c3c */;
            3856: data_o = 32'h00000000 /* 0x3c40 */;
            3857: data_o = 32'h00000000 /* 0x3c44 */;
            3858: data_o = 32'h00000000 /* 0x3c48 */;
            3859: data_o = 32'h00000000 /* 0x3c4c */;
            3860: data_o = 32'h00000000 /* 0x3c50 */;
            3861: data_o = 32'h00000000 /* 0x3c54 */;
            3862: data_o = 32'h00000000 /* 0x3c58 */;
            3863: data_o = 32'h00000000 /* 0x3c5c */;
            3864: data_o = 32'h00000000 /* 0x3c60 */;
            3865: data_o = 32'h00000000 /* 0x3c64 */;
            3866: data_o = 32'h00000000 /* 0x3c68 */;
            3867: data_o = 32'h00000000 /* 0x3c6c */;
            3868: data_o = 32'h00000000 /* 0x3c70 */;
            3869: data_o = 32'h00000000 /* 0x3c74 */;
            3870: data_o = 32'h00000000 /* 0x3c78 */;
            3871: data_o = 32'h00000000 /* 0x3c7c */;
            3872: data_o = 32'h00000000 /* 0x3c80 */;
            3873: data_o = 32'h00000000 /* 0x3c84 */;
            3874: data_o = 32'h00000000 /* 0x3c88 */;
            3875: data_o = 32'h00000000 /* 0x3c8c */;
            3876: data_o = 32'h00000000 /* 0x3c90 */;
            3877: data_o = 32'h00000000 /* 0x3c94 */;
            3878: data_o = 32'h00000000 /* 0x3c98 */;
            3879: data_o = 32'h00000000 /* 0x3c9c */;
            3880: data_o = 32'h00000000 /* 0x3ca0 */;
            3881: data_o = 32'h00000000 /* 0x3ca4 */;
            3882: data_o = 32'h00000000 /* 0x3ca8 */;
            3883: data_o = 32'h00000000 /* 0x3cac */;
            3884: data_o = 32'h00000000 /* 0x3cb0 */;
            3885: data_o = 32'h00000000 /* 0x3cb4 */;
            3886: data_o = 32'h00000000 /* 0x3cb8 */;
            3887: data_o = 32'h00000000 /* 0x3cbc */;
            3888: data_o = 32'h00000000 /* 0x3cc0 */;
            3889: data_o = 32'h00000000 /* 0x3cc4 */;
            3890: data_o = 32'h00000000 /* 0x3cc8 */;
            3891: data_o = 32'h00000000 /* 0x3ccc */;
            3892: data_o = 32'h00000000 /* 0x3cd0 */;
            3893: data_o = 32'h00000000 /* 0x3cd4 */;
            3894: data_o = 32'h00000000 /* 0x3cd8 */;
            3895: data_o = 32'h00000000 /* 0x3cdc */;
            3896: data_o = 32'h00000000 /* 0x3ce0 */;
            3897: data_o = 32'h00000000 /* 0x3ce4 */;
            3898: data_o = 32'h00000000 /* 0x3ce8 */;
            3899: data_o = 32'h00000000 /* 0x3cec */;
            3900: data_o = 32'h00000000 /* 0x3cf0 */;
            3901: data_o = 32'h00000000 /* 0x3cf4 */;
            3902: data_o = 32'h00000000 /* 0x3cf8 */;
            3903: data_o = 32'h00000000 /* 0x3cfc */;
            3904: data_o = 32'h00000000 /* 0x3d00 */;
            3905: data_o = 32'h00000000 /* 0x3d04 */;
            3906: data_o = 32'h00000000 /* 0x3d08 */;
            3907: data_o = 32'h00000000 /* 0x3d0c */;
            3908: data_o = 32'h00000000 /* 0x3d10 */;
            3909: data_o = 32'h00000000 /* 0x3d14 */;
            3910: data_o = 32'h00000000 /* 0x3d18 */;
            3911: data_o = 32'h00000000 /* 0x3d1c */;
            3912: data_o = 32'h00000000 /* 0x3d20 */;
            3913: data_o = 32'h00000000 /* 0x3d24 */;
            3914: data_o = 32'h00000000 /* 0x3d28 */;
            3915: data_o = 32'h00000000 /* 0x3d2c */;
            3916: data_o = 32'h00000000 /* 0x3d30 */;
            3917: data_o = 32'h00000000 /* 0x3d34 */;
            3918: data_o = 32'h00000000 /* 0x3d38 */;
            3919: data_o = 32'h00000000 /* 0x3d3c */;
            3920: data_o = 32'h00000000 /* 0x3d40 */;
            3921: data_o = 32'h00000000 /* 0x3d44 */;
            3922: data_o = 32'h00000000 /* 0x3d48 */;
            3923: data_o = 32'h00000000 /* 0x3d4c */;
            3924: data_o = 32'h00000000 /* 0x3d50 */;
            3925: data_o = 32'h00000000 /* 0x3d54 */;
            3926: data_o = 32'h00000000 /* 0x3d58 */;
            3927: data_o = 32'h00000000 /* 0x3d5c */;
            3928: data_o = 32'h00000000 /* 0x3d60 */;
            3929: data_o = 32'h00000000 /* 0x3d64 */;
            3930: data_o = 32'h00000000 /* 0x3d68 */;
            3931: data_o = 32'h00000000 /* 0x3d6c */;
            3932: data_o = 32'h00000000 /* 0x3d70 */;
            3933: data_o = 32'h00000000 /* 0x3d74 */;
            3934: data_o = 32'h00000000 /* 0x3d78 */;
            3935: data_o = 32'h00000000 /* 0x3d7c */;
            3936: data_o = 32'h00000000 /* 0x3d80 */;
            3937: data_o = 32'h00000000 /* 0x3d84 */;
            3938: data_o = 32'h00000000 /* 0x3d88 */;
            3939: data_o = 32'h00000000 /* 0x3d8c */;
            3940: data_o = 32'h00000000 /* 0x3d90 */;
            3941: data_o = 32'h00000000 /* 0x3d94 */;
            3942: data_o = 32'h00000000 /* 0x3d98 */;
            3943: data_o = 32'h00000000 /* 0x3d9c */;
            3944: data_o = 32'h00000000 /* 0x3da0 */;
            3945: data_o = 32'h00000000 /* 0x3da4 */;
            3946: data_o = 32'h00000000 /* 0x3da8 */;
            3947: data_o = 32'h00000000 /* 0x3dac */;
            3948: data_o = 32'h00000000 /* 0x3db0 */;
            3949: data_o = 32'h00000000 /* 0x3db4 */;
            3950: data_o = 32'h00000000 /* 0x3db8 */;
            3951: data_o = 32'h00000000 /* 0x3dbc */;
            3952: data_o = 32'h00000000 /* 0x3dc0 */;
            3953: data_o = 32'h00000000 /* 0x3dc4 */;
            3954: data_o = 32'h00000000 /* 0x3dc8 */;
            3955: data_o = 32'h00000000 /* 0x3dcc */;
            3956: data_o = 32'h00000000 /* 0x3dd0 */;
            3957: data_o = 32'h00000000 /* 0x3dd4 */;
            3958: data_o = 32'h00000000 /* 0x3dd8 */;
            3959: data_o = 32'h00000000 /* 0x3ddc */;
            3960: data_o = 32'h00000000 /* 0x3de0 */;
            3961: data_o = 32'h00000000 /* 0x3de4 */;
            3962: data_o = 32'h00000000 /* 0x3de8 */;
            3963: data_o = 32'h00000000 /* 0x3dec */;
            3964: data_o = 32'h00000000 /* 0x3df0 */;
            3965: data_o = 32'h00000000 /* 0x3df4 */;
            3966: data_o = 32'h00000000 /* 0x3df8 */;
            3967: data_o = 32'h00000000 /* 0x3dfc */;
            3968: data_o = 32'h00000000 /* 0x3e00 */;
            3969: data_o = 32'h00000000 /* 0x3e04 */;
            3970: data_o = 32'h00000000 /* 0x3e08 */;
            3971: data_o = 32'h00000000 /* 0x3e0c */;
            3972: data_o = 32'h00000000 /* 0x3e10 */;
            3973: data_o = 32'h00000000 /* 0x3e14 */;
            3974: data_o = 32'h00000000 /* 0x3e18 */;
            3975: data_o = 32'h00000000 /* 0x3e1c */;
            3976: data_o = 32'h00000000 /* 0x3e20 */;
            3977: data_o = 32'h00000000 /* 0x3e24 */;
            3978: data_o = 32'h00000000 /* 0x3e28 */;
            3979: data_o = 32'h00000000 /* 0x3e2c */;
            3980: data_o = 32'h00000000 /* 0x3e30 */;
            3981: data_o = 32'h00000000 /* 0x3e34 */;
            3982: data_o = 32'h00000000 /* 0x3e38 */;
            3983: data_o = 32'h00000000 /* 0x3e3c */;
            3984: data_o = 32'h00000000 /* 0x3e40 */;
            3985: data_o = 32'h00000000 /* 0x3e44 */;
            3986: data_o = 32'h00000000 /* 0x3e48 */;
            3987: data_o = 32'h00000000 /* 0x3e4c */;
            3988: data_o = 32'h00000000 /* 0x3e50 */;
            3989: data_o = 32'h00000000 /* 0x3e54 */;
            3990: data_o = 32'h00000000 /* 0x3e58 */;
            3991: data_o = 32'h00000000 /* 0x3e5c */;
            3992: data_o = 32'h00000000 /* 0x3e60 */;
            3993: data_o = 32'h00000000 /* 0x3e64 */;
            3994: data_o = 32'h00000000 /* 0x3e68 */;
            3995: data_o = 32'h00000000 /* 0x3e6c */;
            3996: data_o = 32'h00000000 /* 0x3e70 */;
            3997: data_o = 32'h00000000 /* 0x3e74 */;
            3998: data_o = 32'h00000000 /* 0x3e78 */;
            3999: data_o = 32'h00000000 /* 0x3e7c */;
            4000: data_o = 32'h00000000 /* 0x3e80 */;
            4001: data_o = 32'h00000000 /* 0x3e84 */;
            4002: data_o = 32'h00000000 /* 0x3e88 */;
            4003: data_o = 32'h00000000 /* 0x3e8c */;
            4004: data_o = 32'h00000000 /* 0x3e90 */;
            4005: data_o = 32'h00000000 /* 0x3e94 */;
            4006: data_o = 32'h00000000 /* 0x3e98 */;
            4007: data_o = 32'h00000000 /* 0x3e9c */;
            4008: data_o = 32'h00000000 /* 0x3ea0 */;
            4009: data_o = 32'h00000000 /* 0x3ea4 */;
            4010: data_o = 32'h00000000 /* 0x3ea8 */;
            4011: data_o = 32'h00000000 /* 0x3eac */;
            4012: data_o = 32'h00000000 /* 0x3eb0 */;
            4013: data_o = 32'h00000000 /* 0x3eb4 */;
            4014: data_o = 32'h00000000 /* 0x3eb8 */;
            4015: data_o = 32'h00000000 /* 0x3ebc */;
            4016: data_o = 32'h00000000 /* 0x3ec0 */;
            4017: data_o = 32'h00000000 /* 0x3ec4 */;
            4018: data_o = 32'h00000000 /* 0x3ec8 */;
            4019: data_o = 32'h00000000 /* 0x3ecc */;
            4020: data_o = 32'h00000000 /* 0x3ed0 */;
            4021: data_o = 32'h00000000 /* 0x3ed4 */;
            4022: data_o = 32'h00000000 /* 0x3ed8 */;
            4023: data_o = 32'h00000000 /* 0x3edc */;
            4024: data_o = 32'h00000000 /* 0x3ee0 */;
            4025: data_o = 32'h00000000 /* 0x3ee4 */;
            4026: data_o = 32'h00000000 /* 0x3ee8 */;
            4027: data_o = 32'h00000000 /* 0x3eec */;
            4028: data_o = 32'h00000000 /* 0x3ef0 */;
            4029: data_o = 32'h00000000 /* 0x3ef4 */;
            4030: data_o = 32'h00000000 /* 0x3ef8 */;
            4031: data_o = 32'h00000000 /* 0x3efc */;
            4032: data_o = 32'h00000000 /* 0x3f00 */;
            4033: data_o = 32'h00000000 /* 0x3f04 */;
            4034: data_o = 32'h00000000 /* 0x3f08 */;
            4035: data_o = 32'h00000000 /* 0x3f0c */;
            4036: data_o = 32'h00000000 /* 0x3f10 */;
            4037: data_o = 32'h00000000 /* 0x3f14 */;
            4038: data_o = 32'h00000000 /* 0x3f18 */;
            4039: data_o = 32'h00000000 /* 0x3f1c */;
            4040: data_o = 32'h00000000 /* 0x3f20 */;
            4041: data_o = 32'h00000000 /* 0x3f24 */;
            4042: data_o = 32'h00000000 /* 0x3f28 */;
            4043: data_o = 32'h00000000 /* 0x3f2c */;
            4044: data_o = 32'h00000000 /* 0x3f30 */;
            4045: data_o = 32'h00000000 /* 0x3f34 */;
            4046: data_o = 32'h00000000 /* 0x3f38 */;
            4047: data_o = 32'h00000000 /* 0x3f3c */;
            4048: data_o = 32'h00000000 /* 0x3f40 */;
            4049: data_o = 32'h00000000 /* 0x3f44 */;
            4050: data_o = 32'h00000000 /* 0x3f48 */;
            4051: data_o = 32'h00000000 /* 0x3f4c */;
            4052: data_o = 32'h00000000 /* 0x3f50 */;
            4053: data_o = 32'h00000000 /* 0x3f54 */;
            4054: data_o = 32'h00000000 /* 0x3f58 */;
            4055: data_o = 32'h00000000 /* 0x3f5c */;
            4056: data_o = 32'h00000000 /* 0x3f60 */;
            4057: data_o = 32'h00000000 /* 0x3f64 */;
            4058: data_o = 32'h00000000 /* 0x3f68 */;
            4059: data_o = 32'h00000000 /* 0x3f6c */;
            4060: data_o = 32'h00000000 /* 0x3f70 */;
            4061: data_o = 32'h00000000 /* 0x3f74 */;
            4062: data_o = 32'h00000000 /* 0x3f78 */;
            4063: data_o = 32'h00000000 /* 0x3f7c */;
            4064: data_o = 32'h00000000 /* 0x3f80 */;
            4065: data_o = 32'h00000000 /* 0x3f84 */;
            4066: data_o = 32'h00000000 /* 0x3f88 */;
            4067: data_o = 32'h00000000 /* 0x3f8c */;
            4068: data_o = 32'h00000000 /* 0x3f90 */;
            4069: data_o = 32'h00000000 /* 0x3f94 */;
            4070: data_o = 32'h00000000 /* 0x3f98 */;
            4071: data_o = 32'h00000000 /* 0x3f9c */;
            4072: data_o = 32'h00000000 /* 0x3fa0 */;
            4073: data_o = 32'h00000000 /* 0x3fa4 */;
            4074: data_o = 32'h00000000 /* 0x3fa8 */;
            4075: data_o = 32'h00000000 /* 0x3fac */;
            4076: data_o = 32'h00000000 /* 0x3fb0 */;
            4077: data_o = 32'h00000000 /* 0x3fb4 */;
            4078: data_o = 32'h00000000 /* 0x3fb8 */;
            4079: data_o = 32'h00000000 /* 0x3fbc */;
            4080: data_o = 32'h00000000 /* 0x3fc0 */;
            4081: data_o = 32'h00000000 /* 0x3fc4 */;
            4082: data_o = 32'h00000000 /* 0x3fc8 */;
            4083: data_o = 32'h00000000 /* 0x3fcc */;
            4084: data_o = 32'h00000000 /* 0x3fd0 */;
            4085: data_o = 32'h00000000 /* 0x3fd4 */;
            4086: data_o = 32'h00000000 /* 0x3fd8 */;
            4087: data_o = 32'h00000000 /* 0x3fdc */;
            4088: data_o = 32'h00000000 /* 0x3fe0 */;
            4089: data_o = 32'h00000000 /* 0x3fe4 */;
            4090: data_o = 32'h00000000 /* 0x3fe8 */;
            4091: data_o = 32'h00000000 /* 0x3fec */;
            4092: data_o = 32'h00000000 /* 0x3ff0 */;
            4093: data_o = 32'h00000000 /* 0x3ff4 */;
            4094: data_o = 32'h00000000 /* 0x3ff8 */;
            4095: data_o = 32'h00000000 /* 0x3ffc */;
            default: data_o = '0;
        endcase
    end

endmodule
